module top( n5 , n6 , n15 , n59 , n69 , n72 , n84 , n90 , n97 , 
n107 , n117 , n118 , n124 , n132 , n138 , n152 , n154 , n159 , n182 , 
n187 , n238 , n256 , n269 , n283 , n297 , n317 , n318 , n320 , n323 , 
n328 , n348 , n350 , n357 , n397 , n401 , n445 , n448 , n503 , n508 , 
n527 , n534 , n536 , n550 , n554 , n561 , n587 , n589 , n600 , n614 , 
n618 , n620 , n621 , n624 , n626 , n627 , n632 , n664 , n671 , n677 , 
n684 , n695 , n718 , n720 , n749 , n757 , n763 , n775 , n793 , n795 , 
n814 , n822 , n823 , n824 , n836 , n862 , n865 , n869 , n875 , n884 , 
n891 , n899 , n927 , n928 , n951 , n961 , n982 , n1008 , n1020 , n1024 , 
n1039 , n1057 , n1065 , n1079 , n1095 , n1112 , n1167 , n1177 , n1195 , n1220 , 
n1226 , n1258 , n1268 , n1285 , n1292 , n1309 , n1346 , n1377 , n1382 , n1404 , 
n1406 , n1413 , n1445 , n1447 , n1489 , n1491 , n1500 , n1502 , n1518 , n1519 , 
n1571 , n1574 , n1616 , n1635 , n1638 , n1646 , n1660 , n1669 , n1670 , n1681 , 
n1692 , n1720 , n1742 , n1744 , n1761 , n1785 , n1808 , n1811 , n1819 , n1848 , 
n1849 , n1856 , n1881 , n1888 , n1896 , n1901 , n1906 , n1908 , n1917 , n1918 , 
n1923 , n1932 , n1933 , n1935 , n1980 , n1987 , n1995 , n1997 , n2001 , n2012 , 
n2034 , n2053 , n2056 , n2074 , n2088 , n2113 , n2141 , n2147 , n2150 , n2156 , 
n2159 , n2165 , n2173 , n2192 , n2202 , n2231 , n2245 , n2253 , n2269 , n2303 , 
n2348 , n2382 , n2392 , n2393 , n2422 , n2444 , n2447 , n2467 , n2483 , n2494 , 
n2526 , n2549 , n2552 , n2563 , n2569 , n2610 , n2614 , n2626 , n2629 , n2652 , 
n2665 , n2680 , n2691 , n2703 , n2711 , n2730 , n2798 , n2804 , n2824 , n2825 , 
n2829 , n2846 , n2847 , n2862 , n2873 , n2878 , n2883 , n2884 , n2898 , n2924 , 
n2925 , n2934 , n2939 , n2963 , n3036 , n3048 , n3076 , n3080 , n3084 , n3089 , 
n3105 , n3106 , n3108 , n3131 , n3139 , n3153 , n3163 , n3166 , n3179 , n3185 , 
n3202 , n3214 , n3228 , n3241 , n3259 , n3268 , n3270 , n3281 , n3282 , n3289 , 
n3297 , n3307 , n3312 , n3314 , n3323 , n3345 , n3390 , n3394 , n3425 , n3432 , 
n3433 , n3440 , n3446 , n3460 , n3469 , n3485 , n3515 , n3523 , n3526 , n3553 , 
n3557 , n3573 , n3591 , n3599 , n3612 , n3614 , n3620 , n3624 , n3641 , n3646 , 
n3686 , n3688 , n3717 , n3722 , n3733 , n3755 , n3765 , n3769 , n3772 , n3778 , 
n3782 , n3803 , n3810 , n3822 , n3828 , n3837 , n3858 , n3863 , n3888 , n3907 , 
n3917 , n3928 , n3935 , n3937 , n3942 , n3947 , n3981 , n3993 , n3994 , n3995 , 
n3996 , n4000 , n4015 , n4034 , n4051 , n4054 , n4069 , n4073 , n4077 , n4095 , 
n4130 , n4190 , n4193 , n4213 , n4215 , n4228 , n4257 , n4270 , n4278 , n4300 , 
n4313 , n4317 , n4335 , n4342 , n4350 , n4358 , n4388 , n4393 , n4419 , n4422 , 
n4482 , n4487 , n4515 , n4521 , n4530 , n4554 , n4569 , n4597 , n4611 , n4620 , 
n4622 , n4625 , n4642 , n4647 , n4662 , n4675 , n4708 , n4719 , n4727 , n4733 , 
n4736 , n4743 , n4773 , n4783 , n4805 , n4810 , n4819 , n4836 , n4844 , n4847 , 
n4899 , n4920 , n4924 , n4933 , n4956 , n4958 , n4959 , n5003 , n5008 , n5022 , 
n5024 , n5054 , n5069 , n5088 , n5095 , n5149 , n5150 , n5164 , n5201 , n5211 , 
n5212 , n5226 , n5232 , n5244 , n5251 , n5267 , n5295 , n5299 , n5300 , n5313 , 
n5340 , n5341 , n5360 , n5371 , n5377 , n5385 , n5387 , n5388 , n5442 , n5481 , 
n5510 , n5579 , n5581 , n5593 , n5633 , n5636 , n5638 , n5640 , n5643 , n5649 , 
n5655 , n5661 , n5668 , n5670 , n5685 , n5721 , n5727 , n5732 , n5737 , n5760 , 
n5783 , n5792 , n5831 , n5873 , n5886 , n5888 , n5903 , n5907 , n5922 , n5937 , 
n5941 , n5948 , n5957 , n6036 , n6039 , n6054 , n6074 , n6080 , n6089 , n6105 , 
n6114 , n6127 , n6133 , n6141 , n6145 , n6172 , n6174 , n6196 , n6200 , n6223 , 
n6249 , n6256 , n6259 , n6295 , n6298 , n6306 , n6313 , n6331 , n6334 , n6337 , 
n6349 , n6362 , n6366 , n6390 , n6403 , n6409 , n6427 , n6430 , n6431 , n6440 , 
n6442 , n6451 , n6458 , n6462 , n6470 , n6504 , n6505 , n6526 , n6527 , n6534 , 
n6544 , n6546 , n6555 , n6602 , n6603 , n6626 , n6632 , n6651 , n6687 , n6711 , 
n6734 , n6743 , n6794 , n6803 , n6809 , n6813 , n6815 , n6862 , n6874 , n6888 , 
n6893 , n6919 , n6940 , n6946 , n6957 , n6986 , n7009 , n7014 , n7023 , n7024 , 
n7043 , n7046 , n7047 , n7075 , n7076 , n7094 , n7125 , n7148 , n7150 , n7155 , 
n7180 , n7183 , n7184 , n7209 , n7210 , n7231 , n7241 , n7255 , n7265 , n7267 , 
n7288 , n7314 , n7315 , n7346 , n7354 , n7363 , n7371 , n7386 , n7411 , n7414 , 
n7425 , n7428 , n7434 , n7447 , n7465 , n7473 , n7478 , n7485 , n7502 , n7540 , 
n7553 , n7593 , n7651 , n7655 , n7668 , n7692 , n7701 , n7705 , n7707 , n7708 , 
n7728 , n7735 , n7760 , n7761 , n7787 , n7795 , n7828 , n7852 , n7862 , n7878 , 
n7890 , n7948 , n7987 , n8005 , n8014 , n8030 , n8042 , n8063 , n8067 , n8076 , 
n8095 , n8097 , n8104 , n8109 , n8125 , n8180 , n8183 , n8194 , n8235 , n8242 , 
n8260 , n8264 , n8270 , n8296 , n8297 , n8301 , n8307 , n8314 , n8319 , n8320 , 
n8321 , n8323 , n8365 , n8379 , n8380 , n8384 , n8406 , n8407 , n8430 , n8460 , 
n8485 , n8513 , n8561 , n8566 , n8570 , n8584 , n8606 , n8620 , n8621 , n8628 , 
n8631 , n8685 , n8689 , n8706 , n8713 , n8714 , n8737 , n8771 , n8784 , n8804 , 
n8808 , n8820 , n8834 , n8836 , n8867 , n8873 , n8876 , n8902 , n8919 , n8949 , 
n8958 , n8986 , n8988 , n9011 , n9036 , n9043 , n9067 , n9099 , n9105 , n9115 , 
n9116 , n9132 , n9144 , n9145 , n9163 , n9209 , n9223 , n9228 , n9234 , n9239 , 
n9246 , n9258 , n9274 , n9277 , n9303 , n9310 , n9318 , n9321 , n9336 , n9338 , 
n9358 , n9414 , n9424 , n9469 , n9497 , n9509 , n9517 , n9519 , n9526 , n9532 , 
n9535 , n9554 , n9563 , n9591 , n9593 , n9604 , n9608 , n9619 , n9632 , n9643 , 
n9647 , n9653 , n9655 , n9656 , n9691 , n9708 , n9744 , n9785 , n9796 , n9831 , 
n9835 , n9854 , n9880 , n9898 , n9908 , n9918 , n9929 , n9935 , n9939 , n9945 , 
n9948 , n9959 , n9980 , n9984 , n9985 , n10004 , n10024 , n10034 , n10071 , n10077 , 
n10095 , n10114 , n10117 , n10127 , n10128 , n10139 , n10140 , n10156 , n10158 , n10171 , 
n10172 , n10174 , n10176 , n10193 , n10209 , n10226 , n10251 , n10254 , n10263 , n10269 , 
n10292 , n10296 , n10306 , n10320 , n10327 , n10334 , n10335 , n10352 , n10353 , n10358 , 
n10363 , n10365 , n10393 , n10408 , n10413 , n10417 , n10433 , n10438 , n10451 , n10461 , 
n10471 , n10474 , n10475 , n10477 , n10490 , n10521 , n10551 , n10553 , n10583 , n10615 , 
n10619 , n10620 , n10640 , n10643 , n10676 , n10690 , n10692 , n10728 , n10737 , n10753 , 
n10795 , n10800 , n10825 , n10865 , n10866 , n10868 , n10910 , n10914 , n10949 , n10956 , 
n10966 , n10977 , n10981 , n10990 , n10996 , n11023 , n11031 , n11051 , n11060 , n11062 , 
n11065 , n11132 , n11140 , n11197 , n11208 , n11218 , n11223 , n11227 , n11245 , n11253 , 
n11262 , n11269 , n11328 , n11338 , n11353 , n11360 , n11361 , n11368 , n11373 , n11401 , 
n11407 , n11433 , n11462 , n11485 , n11547 , n11574 , n11585 , n11599 , n11601 , n11610 , 
n11613 , n11614 , n11634 , n11643 , n11653 , n11658 , n11682 , n11685 , n11692 , n11711 , 
n11714 , n11722 , n11736 , n11771 , n11789 , n11792 , n11812 , n11814 , n11839 , n11840 , 
n11847 , n11866 , n11884 , n11886 , n11905 , n11907 , n11963 , n11984 , n11997 , n12024 , 
n12030 , n12032 , n12035 , n12038 , n12049 , n12055 , n12072 , n12105 , n12126 , n12127 , 
n12135 , n12143 , n12165 , n12181 , n12194 , n12196 , n12207 , n12210 , n12220 , n12231 , 
n12242 , n12243 , n12245 , n12259 , n12265 , n12271 , n12312 , n12364 , n12374 , n12380 , 
n12398 , n12399 , n12404 , n12409 , n12426 , n12438 , n12454 , n12464 , n12478 , n12495 , 
n12514 , n12530 , n12561 , n12566 , n12572 , n12587 , n12605 , n12607 , n12625 , n12627 , 
n12638 , n12653 , n12668 , n12669 , n12678 , n12681 , n12686 , n12695 , n12704 , n12707 , 
n12712 , n12713 , n12726 , n12734 , n12737 , n12777 , n12803 , n12805 , n12806 , n12814 , 
n12838 , n12839 , n12870 , n12920 , n12942 , n12946 , n12975 , n12998 , n13004 , n13021 , 
n13048 , n13064 , n13104 , n13114 , n13137 , n13145 , n13161 , n13179 , n13181 , n13210 , 
n13211 , n13215 , n13219 , n13234 , n13235 , n13237 , n13271 , n13276 , n13280 , n13289 , 
n13308 , n13344 , n13345 , n13358 , n13360 , n13364 , n13365 , n13374 , n13380 , n13385 , 
n13389 , n13399 , n13406 , n13410 , n13437 , n13450 , n13453 , n13454 , n13494 , n13504 , 
n13514 , n13526 , n13545 , n13556 , n13559 , n13562 , n13577 , n13604 , n13619 , n13635 , 
n13640 , n13653 , n13654 , n13661 , n13667 , n13679 , n13700 , n13701 , n13725 , n13751 , 
n13800 , n13808 , n13811 , n13833 , n13842 , n13850 , n13859 , n13861 , n13867 , n13910 , 
n13914 , n13932 , n13957 , n13964 , n13975 , n13980 , n13984 , n14008 , n14012 , n14016 , 
n14034 , n14035 , n14040 , n14049 , n14054 , n14073 , n14106 , n14110 , n14112 , n14121 , 
n14131 , n14136 , n14137 , n14166 , n14167 , n14200 , n14212 , n14227 , n14259 , n14262 , 
n14290 , n14311 , n14324 , n14344 , n14348 , n14356 , n14361 , n14363 , n14397 , n14409 , 
n14418 , n14435 , n14477 , n14489 , n14490 , n14503 , n14504 , n14519 , n14520 , n14530 , 
n14555 , n14565 , n14571 , n14584 , n14593 , n14603 , n14613 , n14624 , n14638 , n14655 , 
n14665 , n14670 , n14690 , n14699 , n14711 , n14716 , n14753 , n14777 , n14792 , n14795 , 
n14822 , n14826 , n14828 , n14837 , n14872 , n14880 , n14883 , n14907 , n14925 , n14928 , 
n14934 , n14941 , n14954 , n14958 , n14962 , n14967 , n14985 , n14989 , n14992 , n15007 , 
n15009 , n15010 , n15026 , n15049 , n15059 , n15085 , n15100 , n15115 , n15133 , n15143 , 
n15148 , n15155 , n15164 , n15165 , n15167 , n15178 , n15191 , n15219 , n15231 , n15257 , 
n15271 , n15278 , n15318 , n15338 , n15342 , n15351 , n15363 , n15379 , n15382 , n15396 , 
n15406 , n15409 , n15413 , n15416 , n15434 , n15436 , n15471 , n15484 , n15487 , n15494 , 
n15505 , n15511 , n15534 , n15535 , n15558 , n15580 , n15588 , n15591 , n15592 , n15608 , 
n15609 , n15617 , n15618 , n15650 , n15658 , n15693 , n15694 , n15749 , n15753 , n15758 , 
n15763 , n15787 , n15790 , n15804 , n15815 , n15826 , n15847 , n15855 , n15886 , n15900 , 
n15904 , n15922 , n15937 , n15947 , n15951 , n15986 , n15987 , n15988 , n15993 , n15995 , 
n15999 , n16003 , n16019 , n16024 , n16040 , n16047 , n16070 , n16075 , n16081 , n16091 , 
n16104 , n16113 , n16125 , n16131 , n16132 , n16164 , n16170 , n16187 , n16192 , n16200 , 
n16209 , n16220 , n16223 , n16228 , n16238 , n16239 , n16249 , n16252 , n16275 , n16283 , 
n16285 , n16306 , n16308 , n16324 , n16328 , n16329 , n16334 , n16347 , n16361 , n16382 , 
n16406 , n16411 , n16427 , n16434 , n16441 , n16442 , n16487 , n16500 , n16516 , n16522 , 
n16552 , n16558 , n16562 , n16570 , n16591 , n16601 , n16609 , n16619 , n16623 , n16652 , 
n16656 , n16661 , n16671 , n16676 , n16680 , n16694 , n16703 , n16705 , n16707 , n16708 , 
n16718 , n16737 , n16775 , n16785 , n16789 , n16799 , n16803 , n16815 , n16821 , n16824 , 
n16826 , n16837 , n16852 , n16853 , n16856 , n16873 , n16888 , n16893 , n16900 , n16916 , 
n16927 , n16937 , n16951 , n16986 , n16998 , n17019 , n17028 , n17051 , n17052 , n17055 , 
n17058 , n17068 , n17073 , n17089 , n17109 , n17134 , n17149 , n17156 , n17215 , n17227 , 
n17230 , n17242 , n17255 , n17285 , n17302 , n17305 , n17324 , n17354 , n17368 , n17378 , 
n17388 , n17396 , n17402 , n17417 , n17419 , n17439 , n17444 , n17457 , n17470 , n17471 , 
n17473 , n17495 , n17498 , n17499 , n17509 , n17510 , n17524 , n17527 , n17585 , n17586 , 
n17606 , n17607 , n17617 , n17630 , n17657 , n17673 , n17694 , n17695 , n17712 , n17745 , 
n17768 , n17783 , n17798 , n17808 , n17814 , n17829 , n17843 , n17851 , n17855 , n17867 , 
n17883 , n17910 , n17914 , n17916 , n17943 , n17946 , n17981 , n17995 , n18002 , n18012 , 
n18022 , n18037 , n18087 , n18101 , n18134 , n18156 , n18165 , n18174 , n18203 , n18204 , 
n18207 , n18214 , n18245 , n18253 , n18266 , n18278 , n18292 , n18293 , n18334 , n18376 , 
n18380 , n18388 , n18389 , n18391 , n18394 , n18401 , n18423 , n18435 , n18452 , n18479 , 
n18507 , n18510 , n18516 , n18518 , n18519 , n18534 , n18551 , n18582 , n18590 , n18621 , 
n18627 , n18629 , n18640 , n18645 , n18647 , n18654 , n18667 , n18672 , n18730 , n18792 , 
n18810 , n18812 , n18825 , n18850 , n18903 , n18907 , n18939 , n18955 , n18993 , n19026 , 
n19035 , n19051 , n19066 , n19085 , n19092 , n19095 , n19110 , n19132 , n19146 , n19149 , 
n19202 , n19205 , n19207 , n19211 , n19217 , n19221 , n19229 , n19231 , n19235 , n19238 , 
n19255 , n19261 , n19263 , n19271 , n19274 , n19300 , n19317 , n19356 , n19360 , n19371 , 
n19405 , n19425 , n19452 , n19453 , n19459 , n19477 , n19516 , n19538 , n19542 , n19546 , 
n19572 , n19573 , n19591 , n19592 , n19604 , n19607 , n19615 , n19620 , n19632 , n19648 , 
n19662 , n19671 , n19720 , n19759 , n19776 , n19796 , n19823 , n19880 , n19923 , n19925 , 
n19926 , n19934 , n19943 , n19949 , n19956 , n19980 , n19986 , n20018 , n20032 , n20038 , 
n20041 , n20063 , n20065 , n20080 , n20116 , n20135 , n20155 , n20170 , n20175 , n20181 , 
n20198 , n20210 , n20212 , n20213 , n20231 , n20236 , n20246 , n20262 , n20308 , n20338 , 
n20365 , n20379 , n20390 , n20393 , n20400 , n20410 , n20442 , n20453 , n20466 , n20486 , 
n20495 , n20507 , n20510 , n20545 , n20560 , n20589 , n20593 , n20594 , n20632 , n20664 , 
n20665 , n20673 , n20684 , n20693 , n20727 , n20736 , n20749 , n20753 , n20759 , n20768 , 
n20772 , n20799 , n20800 , n20801 , n20808 , n20812 , n20815 , n20825 , n20827 , n20870 , 
n20881 , n20905 , n20929 , n20931 , n20934 , n20957 , n20976 , n20978 , n20989 , n21013 , 
n21021 , n21064 , n21071 , n21104 , n21122 , n21125 , n21136 , n21177 , n21180 , n21185 , 
n21186 , n21239 , n21261 , n21299 , n21301 , n21313 , n21339 , n21343 , n21356 , n21359 , 
n21362 , n21365 , n21385 , n21389 , n21392 , n21420 , n21421 , n21427 , n21440 , n21444 , 
n21453 , n21455 , n21458 , n21466 , n21470 , n21485 , n21493 , n21508 , n21545 , n21548 , 
n21558 , n21563 , n21569 , n21597 , n21603 , n21615 , n21628 , n21632 , n21653 , n21655 , 
n21686 , n21688 , n21702 , n21706 , n21708 , n21722 , n21756 , n21771 , n21780 , n21787 , 
n21790 , n21801 , n21806 , n21808 , n21813 , n21827 , n21835 , n21862 , n21864 , n21870 , 
n21908 , n21918 , n21960 , n21963 , n21966 , n21970 , n21989 , n22009 , n22040 , n22045 , 
n22075 , n22116 , n22118 , n22121 , n22125 , n22164 , n22167 , n22184 , n22185 , n22205 , 
n22207 , n22218 , n22233 , n22257 , n22270 , n22304 , n22305 , n22316 , n22386 , n22388 , 
n22393 , n22421 , n22422 , n22423 , n22434 , n22443 , n22451 , n22498 , n22512 , n22530 , 
n22541 , n22549 , n22550 , n22564 , n22575 , n22600 , n22603 , n22633 , n22649 , n22665 , 
n22666 , n22667 , n22675 , n22678 , n22701 , n22702 , n22713 , n22715 , n22773 , n22799 , 
n22829 , n22830 , n22845 , n22856 , n22864 , n22866 , n22867 , n22878 , n22886 , n22909 , 
n22913 , n22917 , n22920 , n22922 , n22929 , n22960 , n22962 , n22979 , n22985 , n23023 , 
n23040 , n23043 , n23046 , n23047 , n23052 , n23071 , n23076 , n23097 , n23108 , n23115 , 
n23143 , n23144 , n23145 , n23156 , n23164 , n23165 , n23195 , n23199 , n23204 , n23218 , 
n23232 , n23282 , n23288 , n23304 , n23306 , n23320 , n23326 , n23336 , n23342 , n23374 , 
n23375 , n23400 , n23403 , n23406 , n23407 , n23419 , n23429 , n23431 , n23464 , n23540 , 
n23542 , n23551 , n23558 , n23560 , n23561 , n23565 , n23577 , n23620 , n23643 , n23655 , 
n23681 , n23734 , n23744 , n23749 , n23770 , n23771 , n23787 , n23800 , n23824 , n23832 , 
n23835 , n23838 , n23852 , n23906 , n23922 , n23934 , n23960 , n23997 , n24021 , n24022 , 
n24047 , n24053 , n24056 , n24066 , n24086 , n24100 , n24114 , n24118 , n24132 , n24137 , 
n24144 , n24179 , n24184 , n24213 , n24222 , n24238 , n24246 , n24283 , n24289 , n24304 , 
n24311 , n24338 , n24350 , n24377 , n24398 , n24415 , n24429 , n24455 , n24464 , n24473 , 
n24478 , n24512 , n24515 , n24522 , n24525 , n24526 , n24535 , n24549 , n24569 , n24575 , 
n24578 , n24586 , n24591 , n24628 , n24648 , n24666 , n24687 , n24708 , n24712 , n24744 , 
n24767 , n24770 , n24774 , n24789 , n24794 , n24803 , n24804 , n24807 , n24808 , n24811 , 
n24817 , n24837 , n24841 , n24885 , n24892 , n24895 , n24937 , n24939 , n24946 , n24988 , 
n24999 , n25002 , n25043 , n25089 , n25112 , n25123 , n25171 , n25172 , n25193 , n25235 , 
n25242 , n25251 , n25273 , n25276 , n25291 , n25310 , n25329 , n25334 , n25367 , n25396 , 
n25448 , n25450 , n25487 , n25502 , n25508 , n25509 , n25527 , n25539 , n25559 , n25578 , 
n25585 , n25586 , n25633 , n25641 , n25673 , n25699 , n25716 , n25741 , n25742 , n25758 , 
n25760 , n25764 , n25790 , n25793 , n25805 , n25833 , n25870 , n25889 , n25891 , n25930 , 
n25934 , n25945 , n25952 , n25963 , n25968 , n25989 , n25991 , n26001 , n26002 , n26004 , 
n26007 , n26052 , n26054 , n26072 , n26082 , n26090 , n26094 , n26103 , n26108 , n26114 , 
n26115 , n26121 , n26149 , n26153 , n26155 , n26190 , n26191 , n26197 , n26203 , n26306 , 
n26335 , n26415 , n26425 , n26447 , n26456 , n26466 , n26470 , n26508 , n26526 , n26530 , 
n26541 , n26547 , n26553 , n26571 , n26579 , n26598 , n26636 , n26642 , n26665 , n26670 , 
n26694 , n26700 , n26729 , n26741 , n26747 , n26758 , n26764 , n26778 , n26781 , n26785 , 
n26786 , n26812 , n26837 , n26839 , n26844 , n26863 , n26867 , n26880 , n26885 , n26894 , 
n26908 , n26919 , n26932 , n26940 , n26947 , n26960 , n26961 , n26964 , n26974 , n26996 , 
n27002 , n27034 , n27056 , n27064 , n27070 , n27077 , n27085 , n27090 , n27095 , n27126 , 
n27134 , n27141 , n27160 , n27195 , n27211 , n27223 , n27233 , n27252 , n27254 , n27261 , 
n27305 , n27315 , n27318 , n27322 , n27354 , n27355 , n27356 , n27361 , n27396 , n27410 , 
n27443 , n27453 , n27456 , n27464 , n27467 , n27472 , n27477 , n27492 , n27501 , n27502 , 
n27506 , n27508 , n27524 , n27528 , n27534 , n27547 , n27564 , n27571 , n27572 , n27591 , 
n27601 , n27621 , n27632 , n27636 , n27639 , n27658 , n27713 , n27720 , n27730 , n27736 , 
n27805 , n27829 , n27833 , n27848 , n27882 , n27883 , n27885 , n27895 , n27896 , n27898 , 
n27958 , n27974 , n28006 , n28032 , n28081 , n28098 , n28113 , n28116 , n28124 , n28145 , 
n28146 , n28158 , n28180 , n28188 , n28257 , n28267 , n28278 , n28289 , n28305 , n28320 , 
n28337 , n28340 , n28374 , n28397 , n28399 , n28402 , n28416 , n28417 , n28422 , n28433 , 
n28441 , n28517 , n28537 , n28543 , n28552 , n28562 , n28564 , n28604 , n28606 , n28609 , 
n28613 , n28634 , n28636 , n28638 , n28670 , n28681 , n28703 , n28734 , n28750 , n28754 , 
n28781 , n28783 , n28828 , n28852 , n28856 , n28860 , n28878 , n28943 , n28951 , n28952 , 
n28957 , n28960 , n28983 , n28989 , n29001 , n29023 , n29031 , n29059 , n29070 , n29078 , 
n29090 , n29132 , n29153 , n29182 , n29189 , n29227 , n29229 , n29249 , n29265 , n29293 , 
n29306 , n29314 , n29316 , n29360 , n29369 , n29380 , n29382 , n29390 , n29416 , n29417 , 
n29437 , n29444 , n29447 , n29450 , n29455 , n29470 , n29471 , n29478 , n29547 , n29566 , 
n29569 , n29583 , n29604 , n29615 , n29619 , n29623 , n29650 , n29662 , n29666 , n29667 , 
n29668 , n29677 , n29691 , n29692 , n29702 , n29711 , n29720 , n29763 , n29764 , n29804 , 
n29818 , n29833 , n29838 , n29862 , n29878 , n29883 , n29897 , n29902 , n29933 , n29974 , 
n29988 , n29996 , n30002 , n30009 , n30042 , n30056 , n30067 , n30096 , n30111 , n30150 , 
n30153 , n30158 , n30167 , n30170 , n30172 , n30188 , n30201 , n30245 , n30249 , n30250 , 
n30260 , n30266 , n30269 , n30274 , n30282 , n30287 , n30289 , n30297 , n30318 , n30326 , 
n30343 , n30393 , n30405 , n30411 , n30416 , n30425 , n30432 , n30435 , n30457 , n30458 , 
n30505 , n30514 , n30525 , n30529 , n30534 , n30543 , n30545 , n30562 , n30566 , n30567 , 
n30593 , n30624 , n30625 , n30634 , n30655 , n30664 , n30669 , n30679 , n30685 , n30688 , 
n30706 , n30727 , n30729 , n30769 , n30788 , n30797 , n30798 , n30815 , n30821 , n30831 , 
n30837 , n30845 , n30846 , n30887 , n30892 , n30907 , n30908 , n30925 , n30936 , n30937 , 
n30954 , n30984 , n31012 , n31015 , n31017 , n31019 , n31055 , n31058 , n31060 , n31073 , 
n31077 , n31083 , n31094 , n31108 , n31111 , n31127 , n31134 , n31144 , n31168 , n31181 , 
n31189 , n31194 , n31197 , n31204 , n31217 , n31221 , n31254 , n31264 , n31277 , n31286 , 
n31301 , n31321 , n31326 , n31332 , n31349 , n31351 , n31366 , n31370 , n31373 , n31390 , 
n31396 , n31397 , n31421 , n31426 , n31447 , n31448 , n31466 , n31470 , n31481 , n31484 , 
n31505 , n31534 , n31536 , n31570 , n31591 , n31625 , n31650 , n31686 , n31693 , n31701 , 
n31722 , n31725 , n31727 , n31733 , n31736 , n31741 , n31744 , n31762 , n31763 , n31773 , 
n31783 , n31784 , n31789 , n31824 , n31848 , n31854 , n31889 , n31896 , n31907 , n31910 , 
n31940 , n31945 , n31955 , n31970 , n31981 , n31990 , n32018 , n32023 , n32029 );
    input n15 , n84 , n90 , n97 , n107 , n117 , n124 , n138 , n154 , 
n238 , n256 , n283 , n318 , n320 , n350 , n397 , n445 , n508 , n534 , 
n554 , n561 , n614 , n621 , n624 , n626 , n632 , n664 , n671 , n757 , 
n763 , n775 , n793 , n823 , n862 , n891 , n899 , n1020 , n1039 , n1057 , 
n1095 , n1177 , n1195 , n1285 , n1346 , n1404 , n1518 , n1616 , n1635 , n1669 , 
n1670 , n1692 , n1720 , n1742 , n1819 , n1856 , n1923 , n1935 , n1980 , n1995 , 
n1997 , n2001 , n2150 , n2231 , n2444 , n2447 , n2483 , n2610 , n2629 , n2665 , 
n2798 , n2825 , n2862 , n2883 , n2898 , n2924 , n2925 , n2934 , n2939 , n2963 , 
n3036 , n3076 , n3080 , n3106 , n3108 , n3131 , n3163 , n3166 , n3214 , n3259 , 
n3268 , n3281 , n3289 , n3297 , n3307 , n3312 , n3345 , n3432 , n3440 , n3485 , 
n3515 , n3553 , n3591 , n3599 , n3614 , n3620 , n3641 , n3688 , n3755 , n3765 , 
n3782 , n3810 , n3822 , n3828 , n3837 , n3858 , n3863 , n3907 , n3993 , n3996 , 
n4054 , n4069 , n4130 , n4213 , n4257 , n4278 , n4335 , n4350 , n4358 , n4393 , 
n4554 , n4662 , n4836 , n4844 , n4847 , n4924 , n4956 , n5022 , n5069 , n5149 , 
n5150 , n5251 , n5299 , n5300 , n5313 , n5360 , n5387 , n5388 , n5638 , n5685 , 
n5783 , n5792 , n5831 , n5873 , n5948 , n6036 , n6127 , n6141 , n6145 , n6172 , 
n6196 , n6223 , n6249 , n6256 , n6295 , n6306 , n6331 , n6349 , n6527 , n6534 , 
n6603 , n6626 , n6651 , n6803 , n6874 , n6888 , n6940 , n6957 , n7009 , n7014 , 
n7024 , n7046 , n7180 , n7184 , n7209 , n7210 , n7241 , n7314 , n7315 , n7354 , 
n7414 , n7425 , n7434 , n7447 , n7465 , n7473 , n7593 , n7651 , n7655 , n7692 , 
n7701 , n7705 , n7707 , n7728 , n7760 , n7787 , n7890 , n8005 , n8014 , n8030 , 
n8042 , n8063 , n8097 , n8104 , n8183 , n8260 , n8264 , n8321 , n8407 , n8561 , 
n8584 , n8620 , n8713 , n8714 , n8804 , n8808 , n8834 , n8867 , n8873 , n8919 , 
n8986 , n8988 , n9011 , n9043 , n9116 , n9145 , n9163 , n9209 , n9228 , n9239 , 
n9310 , n9318 , n9321 , n9336 , n9338 , n9358 , n9414 , n9424 , n9469 , n9509 , 
n9591 , n9604 , n9619 , n9653 , n9655 , n9691 , n9744 , n9831 , n9835 , n9935 , 
n9939 , n9948 , n10034 , n10071 , n10114 , n10139 , n10158 , n10269 , n10320 , n10327 , 
n10334 , n10363 , n10393 , n10413 , n10433 , n10451 , n10474 , n10477 , n10490 , n10521 , 
n10619 , n10643 , n10676 , n10737 , n10914 , n10949 , n10981 , n11051 , n11060 , n11065 , 
n11132 , n11140 , n11197 , n11218 , n11223 , n11253 , n11262 , n11360 , n11361 , n11368 , 
n11373 , n11462 , n11574 , n11601 , n11610 , n11643 , n11658 , n11692 , n11711 , n11736 , 
n11771 , n11789 , n11792 , n11847 , n11866 , n11886 , n11905 , n11984 , n12024 , n12030 , 
n12035 , n12055 , n12072 , n12105 , n12143 , n12181 , n12207 , n12210 , n12242 , n12312 , 
n12364 , n12398 , n12399 , n12409 , n12426 , n12478 , n12514 , n12566 , n12605 , n12607 , 
n12625 , n12627 , n12668 , n12712 , n12713 , n12777 , n12803 , n12806 , n12920 , n12946 , 
n12998 , n13137 , n13145 , n13210 , n13271 , n13410 , n13437 , n13454 , n13494 , n13514 , 
n13526 , n13604 , n13635 , n13640 , n13700 , n13701 , n13725 , n13751 , n13800 , n13833 , 
n13859 , n13957 , n13975 , n13980 , n14035 , n14040 , n14106 , n14112 , n14121 , n14136 , 
n14227 , n14290 , n14324 , n14356 , n14361 , n14363 , n14477 , n14489 , n14503 , n14504 , 
n14520 , n14555 , n14624 , n14670 , n14690 , n14711 , n14777 , n14792 , n14795 , n14828 , 
n14872 , n14925 , n14954 , n14962 , n14967 , n14992 , n15009 , n15010 , n15085 , n15100 , 
n15178 , n15191 , n15219 , n15342 , n15363 , n15382 , n15396 , n15413 , n15436 , n15558 , 
n15588 , n15749 , n15758 , n15847 , n15922 , n15987 , n15993 , n15999 , n16019 , n16075 , 
n16113 , n16131 , n16132 , n16200 , n16209 , n16238 , n16283 , n16308 , n16347 , n16406 , 
n16411 , n16441 , n16516 , n16558 , n16570 , n16609 , n16676 , n16785 , n16799 , n16803 , 
n16815 , n16821 , n16856 , n16873 , n16986 , n16998 , n17019 , n17051 , n17068 , n17089 , 
n17109 , n17149 , n17227 , n17255 , n17302 , n17305 , n17368 , n17417 , n17457 , n17499 , 
n17585 , n17617 , n17745 , n17798 , n17843 , n17851 , n17867 , n17910 , n17981 , n17995 , 
n18002 , n18087 , n18165 , n18203 , n18207 , n18253 , n18376 , n18380 , n18388 , n18389 , 
n18391 , n18394 , n18452 , n18507 , n18516 , n18518 , n18534 , n18551 , n18582 , n18645 , 
n18647 , n18667 , n18730 , n18825 , n18850 , n18907 , n18955 , n19035 , n19066 , n19092 , 
n19132 , n19211 , n19217 , n19221 , n19231 , n19238 , n19255 , n19274 , n19300 , n19317 , 
n19356 , n19405 , n19425 , n19516 , n19538 , n19572 , n19592 , n19615 , n19632 , n19720 , 
n19880 , n19943 , n19956 , n20038 , n20041 , n20080 , n20116 , n20135 , n20155 , n20175 , 
n20181 , n20198 , n20210 , n20231 , n20236 , n20262 , n20365 , n20379 , n20390 , n20400 , 
n20442 , n20453 , n20486 , n20495 , n20510 , n20632 , n20664 , n20736 , n20759 , n20799 , 
n20815 , n20825 , n20870 , n20881 , n20905 , n20957 , n20978 , n21064 , n21104 , n21122 , 
n21136 , n21180 , n21185 , n21186 , n21261 , n21301 , n21392 , n21458 , n21466 , n21485 , 
n21493 , n21508 , n21597 , n21603 , n21653 , n21708 , n21771 , n21808 , n21918 , n21960 , 
n21963 , n22045 , n22075 , n22184 , n22233 , n22316 , n22393 , n22421 , n22422 , n22423 , 
n22434 , n22451 , n22512 , n22549 , n22550 , n22665 , n22675 , n22678 , n22845 , n22866 , 
n22867 , n22886 , n22917 , n22922 , n23023 , n23040 , n23043 , n23046 , n23047 , n23052 , 
n23071 , n23097 , n23115 , n23145 , n23195 , n23218 , n23232 , n23306 , n23320 , n23342 , 
n23400 , n23419 , n23561 , n23577 , n23620 , n23643 , n23681 , n23744 , n23770 , n23852 , 
n23934 , n23960 , n24056 , n24066 , n24086 , n24118 , n24132 , n24137 , n24184 , n24213 , 
n24246 , n24289 , n24304 , n24350 , n24377 , n24415 , n24429 , n24455 , n24464 , n24512 , 
n24522 , n24525 , n24569 , n24578 , n24687 , n24712 , n24794 , n24807 , n24837 , n24939 , 
n24988 , n25089 , n25123 , n25242 , n25276 , n25291 , n25334 , n25527 , n25585 , n25699 , 
n25758 , n25760 , n25793 , n25805 , n25889 , n25991 , n26002 , n26004 , n26052 , n26072 , 
n26082 , n26114 , n26115 , n26191 , n26203 , n26306 , n26456 , n26541 , n26598 , n26636 , 
n26665 , n26670 , n26700 , n26758 , n26786 , n26863 , n26867 , n26894 , n26961 , n26974 , 
n26996 , n27002 , n27034 , n27064 , n27077 , n27126 , n27233 , n27318 , n27322 , n27354 , 
n27355 , n27443 , n27453 , n27501 , n27534 , n27591 , n27632 , n27805 , n27829 , n27848 , 
n27883 , n27885 , n27896 , n27974 , n28006 , n28081 , n28113 , n28158 , n28180 , n28267 , 
n28305 , n28397 , n28402 , n28417 , n28433 , n28441 , n28517 , n28562 , n28634 , n28638 , 
n28734 , n28781 , n28828 , n28856 , n28878 , n28951 , n28983 , n29059 , n29090 , n29132 , 
n29153 , n29249 , n29293 , n29380 , n29390 , n29437 , n29444 , n29447 , n29471 , n29569 , 
n29604 , n29615 , n29667 , n29668 , n29702 , n29764 , n29818 , n29878 , n29897 , n29902 , 
n29933 , n29974 , n30002 , n30067 , n30096 , n30158 , n30167 , n30201 , n30245 , n30274 , 
n30287 , n30297 , n30326 , n30343 , n30405 , n30411 , n30425 , n30457 , n30458 , n30505 , 
n30514 , n30525 , n30529 , n30534 , n30562 , n30593 , n30664 , n30669 , n30685 , n30688 , 
n30706 , n30769 , n30831 , n30887 , n30908 , n30936 , n31019 , n31060 , n31094 , n31108 , 
n31111 , n31168 , n31204 , n31301 , n31326 , n31366 , n31426 , n31448 , n31470 , n31481 , 
n31591 , n31722 , n31725 , n31727 , n31773 , n31783 , n31889 , n31896 , n31910 , n31940 , 
n31970 ;
    output n5 , n6 , n59 , n69 , n72 , n118 , n132 , n152 , n159 , 
n182 , n187 , n269 , n297 , n317 , n323 , n328 , n348 , n357 , n401 , 
n448 , n503 , n527 , n536 , n550 , n587 , n589 , n600 , n618 , n620 , 
n627 , n677 , n684 , n695 , n718 , n720 , n749 , n795 , n814 , n822 , 
n824 , n836 , n865 , n869 , n875 , n884 , n927 , n928 , n951 , n961 , 
n982 , n1008 , n1024 , n1065 , n1079 , n1112 , n1167 , n1220 , n1226 , n1258 , 
n1268 , n1292 , n1309 , n1377 , n1382 , n1406 , n1413 , n1445 , n1447 , n1489 , 
n1491 , n1500 , n1502 , n1519 , n1571 , n1574 , n1638 , n1646 , n1660 , n1681 , 
n1744 , n1761 , n1785 , n1808 , n1811 , n1848 , n1849 , n1881 , n1888 , n1896 , 
n1901 , n1906 , n1908 , n1917 , n1918 , n1932 , n1933 , n1987 , n2012 , n2034 , 
n2053 , n2056 , n2074 , n2088 , n2113 , n2141 , n2147 , n2156 , n2159 , n2165 , 
n2173 , n2192 , n2202 , n2245 , n2253 , n2269 , n2303 , n2348 , n2382 , n2392 , 
n2393 , n2422 , n2467 , n2494 , n2526 , n2549 , n2552 , n2563 , n2569 , n2614 , 
n2626 , n2652 , n2680 , n2691 , n2703 , n2711 , n2730 , n2804 , n2824 , n2829 , 
n2846 , n2847 , n2873 , n2878 , n2884 , n3048 , n3084 , n3089 , n3105 , n3139 , 
n3153 , n3179 , n3185 , n3202 , n3228 , n3241 , n3270 , n3282 , n3314 , n3323 , 
n3390 , n3394 , n3425 , n3433 , n3446 , n3460 , n3469 , n3523 , n3526 , n3557 , 
n3573 , n3612 , n3624 , n3646 , n3686 , n3717 , n3722 , n3733 , n3769 , n3772 , 
n3778 , n3803 , n3888 , n3917 , n3928 , n3935 , n3937 , n3942 , n3947 , n3981 , 
n3994 , n3995 , n4000 , n4015 , n4034 , n4051 , n4073 , n4077 , n4095 , n4190 , 
n4193 , n4215 , n4228 , n4270 , n4300 , n4313 , n4317 , n4342 , n4388 , n4419 , 
n4422 , n4482 , n4487 , n4515 , n4521 , n4530 , n4569 , n4597 , n4611 , n4620 , 
n4622 , n4625 , n4642 , n4647 , n4675 , n4708 , n4719 , n4727 , n4733 , n4736 , 
n4743 , n4773 , n4783 , n4805 , n4810 , n4819 , n4899 , n4920 , n4933 , n4958 , 
n4959 , n5003 , n5008 , n5024 , n5054 , n5088 , n5095 , n5164 , n5201 , n5211 , 
n5212 , n5226 , n5232 , n5244 , n5267 , n5295 , n5340 , n5341 , n5371 , n5377 , 
n5385 , n5442 , n5481 , n5510 , n5579 , n5581 , n5593 , n5633 , n5636 , n5640 , 
n5643 , n5649 , n5655 , n5661 , n5668 , n5670 , n5721 , n5727 , n5732 , n5737 , 
n5760 , n5886 , n5888 , n5903 , n5907 , n5922 , n5937 , n5941 , n5957 , n6039 , 
n6054 , n6074 , n6080 , n6089 , n6105 , n6114 , n6133 , n6174 , n6200 , n6259 , 
n6298 , n6313 , n6334 , n6337 , n6362 , n6366 , n6390 , n6403 , n6409 , n6427 , 
n6430 , n6431 , n6440 , n6442 , n6451 , n6458 , n6462 , n6470 , n6504 , n6505 , 
n6526 , n6544 , n6546 , n6555 , n6602 , n6632 , n6687 , n6711 , n6734 , n6743 , 
n6794 , n6809 , n6813 , n6815 , n6862 , n6893 , n6919 , n6946 , n6986 , n7023 , 
n7043 , n7047 , n7075 , n7076 , n7094 , n7125 , n7148 , n7150 , n7155 , n7183 , 
n7231 , n7255 , n7265 , n7267 , n7288 , n7346 , n7363 , n7371 , n7386 , n7411 , 
n7428 , n7478 , n7485 , n7502 , n7540 , n7553 , n7668 , n7708 , n7735 , n7761 , 
n7795 , n7828 , n7852 , n7862 , n7878 , n7948 , n7987 , n8067 , n8076 , n8095 , 
n8109 , n8125 , n8180 , n8194 , n8235 , n8242 , n8270 , n8296 , n8297 , n8301 , 
n8307 , n8314 , n8319 , n8320 , n8323 , n8365 , n8379 , n8380 , n8384 , n8406 , 
n8430 , n8460 , n8485 , n8513 , n8566 , n8570 , n8606 , n8621 , n8628 , n8631 , 
n8685 , n8689 , n8706 , n8737 , n8771 , n8784 , n8820 , n8836 , n8876 , n8902 , 
n8949 , n8958 , n9036 , n9067 , n9099 , n9105 , n9115 , n9132 , n9144 , n9223 , 
n9234 , n9246 , n9258 , n9274 , n9277 , n9303 , n9497 , n9517 , n9519 , n9526 , 
n9532 , n9535 , n9554 , n9563 , n9593 , n9608 , n9632 , n9643 , n9647 , n9656 , 
n9708 , n9785 , n9796 , n9854 , n9880 , n9898 , n9908 , n9918 , n9929 , n9945 , 
n9959 , n9980 , n9984 , n9985 , n10004 , n10024 , n10077 , n10095 , n10117 , n10127 , 
n10128 , n10140 , n10156 , n10171 , n10172 , n10174 , n10176 , n10193 , n10209 , n10226 , 
n10251 , n10254 , n10263 , n10292 , n10296 , n10306 , n10335 , n10352 , n10353 , n10358 , 
n10365 , n10408 , n10417 , n10438 , n10461 , n10471 , n10475 , n10551 , n10553 , n10583 , 
n10615 , n10620 , n10640 , n10690 , n10692 , n10728 , n10753 , n10795 , n10800 , n10825 , 
n10865 , n10866 , n10868 , n10910 , n10956 , n10966 , n10977 , n10990 , n10996 , n11023 , 
n11031 , n11062 , n11208 , n11227 , n11245 , n11269 , n11328 , n11338 , n11353 , n11401 , 
n11407 , n11433 , n11485 , n11547 , n11585 , n11599 , n11613 , n11614 , n11634 , n11653 , 
n11682 , n11685 , n11714 , n11722 , n11812 , n11814 , n11839 , n11840 , n11884 , n11907 , 
n11963 , n11997 , n12032 , n12038 , n12049 , n12126 , n12127 , n12135 , n12165 , n12194 , 
n12196 , n12220 , n12231 , n12243 , n12245 , n12259 , n12265 , n12271 , n12374 , n12380 , 
n12404 , n12438 , n12454 , n12464 , n12495 , n12530 , n12561 , n12572 , n12587 , n12638 , 
n12653 , n12669 , n12678 , n12681 , n12686 , n12695 , n12704 , n12707 , n12726 , n12734 , 
n12737 , n12805 , n12814 , n12838 , n12839 , n12870 , n12942 , n12975 , n13004 , n13021 , 
n13048 , n13064 , n13104 , n13114 , n13161 , n13179 , n13181 , n13211 , n13215 , n13219 , 
n13234 , n13235 , n13237 , n13276 , n13280 , n13289 , n13308 , n13344 , n13345 , n13358 , 
n13360 , n13364 , n13365 , n13374 , n13380 , n13385 , n13389 , n13399 , n13406 , n13450 , 
n13453 , n13504 , n13545 , n13556 , n13559 , n13562 , n13577 , n13619 , n13653 , n13654 , 
n13661 , n13667 , n13679 , n13808 , n13811 , n13842 , n13850 , n13861 , n13867 , n13910 , 
n13914 , n13932 , n13964 , n13984 , n14008 , n14012 , n14016 , n14034 , n14049 , n14054 , 
n14073 , n14110 , n14131 , n14137 , n14166 , n14167 , n14200 , n14212 , n14259 , n14262 , 
n14311 , n14344 , n14348 , n14397 , n14409 , n14418 , n14435 , n14490 , n14519 , n14530 , 
n14565 , n14571 , n14584 , n14593 , n14603 , n14613 , n14638 , n14655 , n14665 , n14699 , 
n14716 , n14753 , n14822 , n14826 , n14837 , n14880 , n14883 , n14907 , n14928 , n14934 , 
n14941 , n14958 , n14985 , n14989 , n15007 , n15026 , n15049 , n15059 , n15115 , n15133 , 
n15143 , n15148 , n15155 , n15164 , n15165 , n15167 , n15231 , n15257 , n15271 , n15278 , 
n15318 , n15338 , n15351 , n15379 , n15406 , n15409 , n15416 , n15434 , n15471 , n15484 , 
n15487 , n15494 , n15505 , n15511 , n15534 , n15535 , n15580 , n15591 , n15592 , n15608 , 
n15609 , n15617 , n15618 , n15650 , n15658 , n15693 , n15694 , n15753 , n15763 , n15787 , 
n15790 , n15804 , n15815 , n15826 , n15855 , n15886 , n15900 , n15904 , n15937 , n15947 , 
n15951 , n15986 , n15988 , n15995 , n16003 , n16024 , n16040 , n16047 , n16070 , n16081 , 
n16091 , n16104 , n16125 , n16164 , n16170 , n16187 , n16192 , n16220 , n16223 , n16228 , 
n16239 , n16249 , n16252 , n16275 , n16285 , n16306 , n16324 , n16328 , n16329 , n16334 , 
n16361 , n16382 , n16427 , n16434 , n16442 , n16487 , n16500 , n16522 , n16552 , n16562 , 
n16591 , n16601 , n16619 , n16623 , n16652 , n16656 , n16661 , n16671 , n16680 , n16694 , 
n16703 , n16705 , n16707 , n16708 , n16718 , n16737 , n16775 , n16789 , n16824 , n16826 , 
n16837 , n16852 , n16853 , n16888 , n16893 , n16900 , n16916 , n16927 , n16937 , n16951 , 
n17028 , n17052 , n17055 , n17058 , n17073 , n17134 , n17156 , n17215 , n17230 , n17242 , 
n17285 , n17324 , n17354 , n17378 , n17388 , n17396 , n17402 , n17419 , n17439 , n17444 , 
n17470 , n17471 , n17473 , n17495 , n17498 , n17509 , n17510 , n17524 , n17527 , n17586 , 
n17606 , n17607 , n17630 , n17657 , n17673 , n17694 , n17695 , n17712 , n17768 , n17783 , 
n17808 , n17814 , n17829 , n17855 , n17883 , n17914 , n17916 , n17943 , n17946 , n18012 , 
n18022 , n18037 , n18101 , n18134 , n18156 , n18174 , n18204 , n18214 , n18245 , n18266 , 
n18278 , n18292 , n18293 , n18334 , n18401 , n18423 , n18435 , n18479 , n18510 , n18519 , 
n18590 , n18621 , n18627 , n18629 , n18640 , n18654 , n18672 , n18792 , n18810 , n18812 , 
n18903 , n18939 , n18993 , n19026 , n19051 , n19085 , n19095 , n19110 , n19146 , n19149 , 
n19202 , n19205 , n19207 , n19229 , n19235 , n19261 , n19263 , n19271 , n19360 , n19371 , 
n19452 , n19453 , n19459 , n19477 , n19542 , n19546 , n19573 , n19591 , n19604 , n19607 , 
n19620 , n19648 , n19662 , n19671 , n19759 , n19776 , n19796 , n19823 , n19923 , n19925 , 
n19926 , n19934 , n19949 , n19980 , n19986 , n20018 , n20032 , n20063 , n20065 , n20170 , 
n20212 , n20213 , n20246 , n20308 , n20338 , n20393 , n20410 , n20466 , n20507 , n20545 , 
n20560 , n20589 , n20593 , n20594 , n20665 , n20673 , n20684 , n20693 , n20727 , n20749 , 
n20753 , n20768 , n20772 , n20800 , n20801 , n20808 , n20812 , n20827 , n20929 , n20931 , 
n20934 , n20976 , n20989 , n21013 , n21021 , n21071 , n21125 , n21177 , n21239 , n21299 , 
n21313 , n21339 , n21343 , n21356 , n21359 , n21362 , n21365 , n21385 , n21389 , n21420 , 
n21421 , n21427 , n21440 , n21444 , n21453 , n21455 , n21470 , n21545 , n21548 , n21558 , 
n21563 , n21569 , n21615 , n21628 , n21632 , n21655 , n21686 , n21688 , n21702 , n21706 , 
n21722 , n21756 , n21780 , n21787 , n21790 , n21801 , n21806 , n21813 , n21827 , n21835 , 
n21862 , n21864 , n21870 , n21908 , n21966 , n21970 , n21989 , n22009 , n22040 , n22116 , 
n22118 , n22121 , n22125 , n22164 , n22167 , n22185 , n22205 , n22207 , n22218 , n22257 , 
n22270 , n22304 , n22305 , n22386 , n22388 , n22443 , n22498 , n22530 , n22541 , n22564 , 
n22575 , n22600 , n22603 , n22633 , n22649 , n22666 , n22667 , n22701 , n22702 , n22713 , 
n22715 , n22773 , n22799 , n22829 , n22830 , n22856 , n22864 , n22878 , n22909 , n22913 , 
n22920 , n22929 , n22960 , n22962 , n22979 , n22985 , n23076 , n23108 , n23143 , n23144 , 
n23156 , n23164 , n23165 , n23199 , n23204 , n23282 , n23288 , n23304 , n23326 , n23336 , 
n23374 , n23375 , n23403 , n23406 , n23407 , n23429 , n23431 , n23464 , n23540 , n23542 , 
n23551 , n23558 , n23560 , n23565 , n23655 , n23734 , n23749 , n23771 , n23787 , n23800 , 
n23824 , n23832 , n23835 , n23838 , n23906 , n23922 , n23997 , n24021 , n24022 , n24047 , 
n24053 , n24100 , n24114 , n24144 , n24179 , n24222 , n24238 , n24283 , n24311 , n24338 , 
n24398 , n24473 , n24478 , n24515 , n24526 , n24535 , n24549 , n24575 , n24586 , n24591 , 
n24628 , n24648 , n24666 , n24708 , n24744 , n24767 , n24770 , n24774 , n24789 , n24803 , 
n24804 , n24808 , n24811 , n24817 , n24841 , n24885 , n24892 , n24895 , n24937 , n24946 , 
n24999 , n25002 , n25043 , n25112 , n25171 , n25172 , n25193 , n25235 , n25251 , n25273 , 
n25310 , n25329 , n25367 , n25396 , n25448 , n25450 , n25487 , n25502 , n25508 , n25509 , 
n25539 , n25559 , n25578 , n25586 , n25633 , n25641 , n25673 , n25716 , n25741 , n25742 , 
n25764 , n25790 , n25833 , n25870 , n25891 , n25930 , n25934 , n25945 , n25952 , n25963 , 
n25968 , n25989 , n26001 , n26007 , n26054 , n26090 , n26094 , n26103 , n26108 , n26121 , 
n26149 , n26153 , n26155 , n26190 , n26197 , n26335 , n26415 , n26425 , n26447 , n26466 , 
n26470 , n26508 , n26526 , n26530 , n26547 , n26553 , n26571 , n26579 , n26642 , n26694 , 
n26729 , n26741 , n26747 , n26764 , n26778 , n26781 , n26785 , n26812 , n26837 , n26839 , 
n26844 , n26880 , n26885 , n26908 , n26919 , n26932 , n26940 , n26947 , n26960 , n26964 , 
n27056 , n27070 , n27085 , n27090 , n27095 , n27134 , n27141 , n27160 , n27195 , n27211 , 
n27223 , n27252 , n27254 , n27261 , n27305 , n27315 , n27356 , n27361 , n27396 , n27410 , 
n27456 , n27464 , n27467 , n27472 , n27477 , n27492 , n27502 , n27506 , n27508 , n27524 , 
n27528 , n27547 , n27564 , n27571 , n27572 , n27601 , n27621 , n27636 , n27639 , n27658 , 
n27713 , n27720 , n27730 , n27736 , n27833 , n27882 , n27895 , n27898 , n27958 , n28032 , 
n28098 , n28116 , n28124 , n28145 , n28146 , n28188 , n28257 , n28278 , n28289 , n28320 , 
n28337 , n28340 , n28374 , n28399 , n28416 , n28422 , n28537 , n28543 , n28552 , n28564 , 
n28604 , n28606 , n28609 , n28613 , n28636 , n28670 , n28681 , n28703 , n28750 , n28754 , 
n28783 , n28852 , n28860 , n28943 , n28952 , n28957 , n28960 , n28989 , n29001 , n29023 , 
n29031 , n29070 , n29078 , n29182 , n29189 , n29227 , n29229 , n29265 , n29306 , n29314 , 
n29316 , n29360 , n29369 , n29382 , n29416 , n29417 , n29450 , n29455 , n29470 , n29478 , 
n29547 , n29566 , n29583 , n29619 , n29623 , n29650 , n29662 , n29666 , n29677 , n29691 , 
n29692 , n29711 , n29720 , n29763 , n29804 , n29833 , n29838 , n29862 , n29883 , n29988 , 
n29996 , n30009 , n30042 , n30056 , n30111 , n30150 , n30153 , n30170 , n30172 , n30188 , 
n30249 , n30250 , n30260 , n30266 , n30269 , n30282 , n30289 , n30318 , n30393 , n30416 , 
n30432 , n30435 , n30543 , n30545 , n30566 , n30567 , n30624 , n30625 , n30634 , n30655 , 
n30679 , n30727 , n30729 , n30788 , n30797 , n30798 , n30815 , n30821 , n30837 , n30845 , 
n30846 , n30892 , n30907 , n30925 , n30937 , n30954 , n30984 , n31012 , n31015 , n31017 , 
n31055 , n31058 , n31073 , n31077 , n31083 , n31127 , n31134 , n31144 , n31181 , n31189 , 
n31194 , n31197 , n31217 , n31221 , n31254 , n31264 , n31277 , n31286 , n31321 , n31332 , 
n31349 , n31351 , n31370 , n31373 , n31390 , n31396 , n31397 , n31421 , n31447 , n31466 , 
n31484 , n31505 , n31534 , n31536 , n31570 , n31625 , n31650 , n31686 , n31693 , n31701 , 
n31733 , n31736 , n31741 , n31744 , n31762 , n31763 , n31784 , n31789 , n31824 , n31848 , 
n31854 , n31907 , n31945 , n31955 , n31981 , n31990 , n32018 , n32023 , n32029 ;
    wire n0 , n1 , n2 , n3 , n4 , n7 , n8 , n9 , n10 , 
n11 , n12 , n13 , n14 , n16 , n17 , n18 , n19 , n20 , n21 , 
n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , 
n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , 
n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , 
n52 , n53 , n54 , n55 , n56 , n57 , n58 , n60 , n61 , n62 , 
n63 , n64 , n65 , n66 , n67 , n68 , n70 , n71 , n73 , n74 , 
n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n85 , 
n86 , n87 , n88 , n89 , n91 , n92 , n93 , n94 , n95 , n96 , 
n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n108 , 
n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n119 , n120 , 
n121 , n122 , n123 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , 
n133 , n134 , n135 , n136 , n137 , n139 , n140 , n141 , n142 , n143 , 
n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n153 , n155 , 
n156 , n157 , n158 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
n177 , n178 , n179 , n180 , n181 , n183 , n184 , n185 , n186 , n188 , 
n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , 
n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , 
n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , 
n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , 
n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n239 , 
n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
n250 , n251 , n252 , n253 , n254 , n255 , n257 , n258 , n259 , n260 , 
n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n270 , n271 , 
n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , 
n282 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
n293 , n294 , n295 , n296 , n298 , n299 , n300 , n301 , n302 , n303 , 
n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , 
n314 , n315 , n316 , n319 , n321 , n322 , n324 , n325 , n326 , n327 , 
n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , 
n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n349 , 
n351 , n352 , n353 , n354 , n355 , n356 , n358 , n359 , n360 , n361 , 
n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , 
n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , 
n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , 
n392 , n393 , n394 , n395 , n396 , n398 , n399 , n400 , n402 , n403 , 
n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , 
n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , 
n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , 
n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , 
n444 , n446 , n447 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , 
n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , 
n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , 
n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , 
n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , 
n496 , n497 , n498 , n499 , n500 , n501 , n502 , n504 , n505 , n506 , 
n507 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , 
n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n528 , 
n529 , n530 , n531 , n532 , n533 , n535 , n537 , n538 , n539 , n540 , 
n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n551 , 
n552 , n553 , n555 , n556 , n557 , n558 , n559 , n560 , n562 , n563 , 
n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , 
n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , 
n584 , n585 , n586 , n588 , n590 , n591 , n592 , n593 , n594 , n595 , 
n596 , n597 , n598 , n599 , n601 , n602 , n603 , n604 , n605 , n606 , 
n607 , n608 , n609 , n610 , n611 , n612 , n613 , n615 , n616 , n617 , 
n619 , n622 , n623 , n625 , n628 , n629 , n630 , n631 , n633 , n634 , 
n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n665 , 
n666 , n667 , n668 , n669 , n670 , n672 , n673 , n674 , n675 , n676 , 
n678 , n679 , n680 , n681 , n682 , n683 , n685 , n686 , n687 , n688 , 
n689 , n690 , n691 , n692 , n693 , n694 , n696 , n697 , n698 , n699 , 
n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n719 , n721 , 
n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , 
n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , 
n742 , n743 , n744 , n745 , n746 , n747 , n748 , n750 , n751 , n752 , 
n753 , n754 , n755 , n756 , n758 , n759 , n760 , n761 , n762 , n764 , 
n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , 
n786 , n787 , n788 , n789 , n790 , n791 , n792 , n794 , n796 , n797 , 
n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , 
n808 , n809 , n810 , n811 , n812 , n813 , n815 , n816 , n817 , n818 , 
n819 , n820 , n821 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , 
n832 , n833 , n834 , n835 , n837 , n838 , n839 , n840 , n841 , n842 , 
n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , 
n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n863 , 
n864 , n866 , n867 , n868 , n870 , n871 , n872 , n873 , n874 , n876 , 
n877 , n878 , n879 , n880 , n881 , n882 , n883 , n885 , n886 , n887 , 
n888 , n889 , n890 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , 
n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
n920 , n921 , n922 , n923 , n924 , n925 , n926 , n929 , n930 , n931 , 
n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , 
n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n952 , 
n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n962 , n963 , 
n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , 
n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n983 , n984 , 
n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , 
n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , 
n1005 , n1006 , n1007 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , 
n1016 , n1017 , n1018 , n1019 , n1021 , n1022 , n1023 , n1025 , n1026 , n1027 , 
n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , 
n1038 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , 
n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1058 , n1059 , 
n1060 , n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 , n1069 , n1070 , 
n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1080 , n1081 , 
n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , 
n1092 , n1093 , n1094 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1113 , 
n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , 
n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , 
n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , 
n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , 
n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , 
n1164 , n1165 , n1166 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , 
n1175 , n1176 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , 
n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1196 , 
n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , 
n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , 
n1217 , n1218 , n1219 , n1221 , n1222 , n1223 , n1224 , n1225 , n1227 , n1228 , 
n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , 
n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1259 , 
n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1269 , n1270 , 
n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
n1281 , n1282 , n1283 , n1284 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , 
n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , 
n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1310 , n1311 , n1312 , n1313 , 
n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , 
n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , 
n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , 
n1344 , n1345 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , 
n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , 
n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , 
n1375 , n1376 , n1378 , n1379 , n1380 , n1381 , n1383 , n1384 , n1385 , n1386 , 
n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , 
n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1405 , n1407 , n1408 , 
n1409 , n1410 , n1411 , n1412 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
n1440 , n1441 , n1442 , n1443 , n1444 , n1446 , n1448 , n1449 , n1450 , n1451 , 
n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , 
n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , 
n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , 
n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1490 , n1492 , n1493 , 
n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1501 , n1503 , n1504 , n1505 , 
n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , 
n1516 , n1517 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , 
n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , 
n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , 
n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , 
n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , 
n1568 , n1569 , n1570 , n1572 , n1573 , n1575 , n1576 , n1577 , n1578 , n1579 , 
n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1617 , n1618 , n1619 , n1620 , 
n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
n1631 , n1632 , n1633 , n1634 , n1636 , n1637 , n1639 , n1640 , n1641 , n1642 , 
n1643 , n1644 , n1645 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , 
n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1661 , n1662 , n1663 , n1664 , 
n1665 , n1666 , n1667 , n1668 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , 
n1677 , n1678 , n1679 , n1680 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , 
n1688 , n1689 , n1690 , n1691 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , 
n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , 
n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
n1719 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
n1740 , n1741 , n1743 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , 
n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1762 , 
n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , 
n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , 
n1783 , n1784 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , 
n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , 
n1804 , n1805 , n1806 , n1807 , n1809 , n1810 , n1812 , n1813 , n1814 , n1815 , 
n1816 , n1817 , n1818 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , 
n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , 
n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , 
n1847 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1857 , n1858 , n1859 , 
n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
n1880 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1889 , n1890 , n1891 , 
n1892 , n1893 , n1894 , n1895 , n1897 , n1898 , n1899 , n1900 , n1902 , n1903 , 
n1904 , n1905 , n1907 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , 
n1916 , n1919 , n1920 , n1921 , n1922 , n1924 , n1925 , n1926 , n1927 , n1928 , 
n1929 , n1930 , n1931 , n1934 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , 
n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , 
n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , 
n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , 
n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1981 , n1982 , 
n1983 , n1984 , n1985 , n1986 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , 
n1994 , n1996 , n1998 , n1999 , n2000 , n2002 , n2003 , n2004 , n2005 , n2006 , 
n2007 , n2008 , n2009 , n2010 , n2011 , n2013 , n2014 , n2015 , n2016 , n2017 , 
n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , 
n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2035 , n2036 , n2037 , n2038 , 
n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , 
n2049 , n2050 , n2051 , n2052 , n2054 , n2055 , n2057 , n2058 , n2059 , n2060 , 
n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
n2071 , n2072 , n2073 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , 
n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2089 , n2090 , n2091 , n2092 , 
n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , 
n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , 
n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , 
n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , 
n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2142 , n2143 , n2144 , 
n2145 , n2146 , n2148 , n2149 , n2151 , n2152 , n2153 , n2154 , n2155 , n2157 , 
n2158 , n2160 , n2161 , n2162 , n2163 , n2164 , n2166 , n2167 , n2168 , n2169 , 
n2170 , n2171 , n2172 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
n2191 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , 
n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , 
n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , 
n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2232 , n2233 , 
n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , 
n2244 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2254 , n2255 , 
n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , 
n2266 , n2267 , n2268 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , 
n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2304 , n2305 , n2306 , n2307 , 
n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , 
n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , 
n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , 
n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , 
n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
n2379 , n2380 , n2381 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
n2390 , n2391 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , 
n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , 
n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , 
n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , 
n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , 
n2443 , n2445 , n2446 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , 
n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , 
n2465 , n2466 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , 
n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2484 , n2485 , n2486 , 
n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2495 , n2496 , n2497 , 
n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , 
n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , 
n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2527 , n2528 , 
n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , 
n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , 
n2550 , n2551 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
n2561 , n2562 , n2564 , n2565 , n2566 , n2567 , n2568 , n2570 , n2571 , n2572 , 
n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , 
n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , 
n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , 
n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2611 , n2612 , n2613 , 
n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , 
n2625 , n2627 , n2628 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
n2647 , n2648 , n2649 , n2650 , n2651 , n2653 , n2654 , n2655 , n2656 , n2657 , 
n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2666 , n2667 , n2668 , 
n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , 
n2679 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
n2690 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
n2701 , n2702 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2712 , 
n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , 
n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2731 , n2732 , n2733 , 
n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , 
n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , 
n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , 
n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , 
n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , 
n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , 
n2794 , n2795 , n2796 , n2797 , n2799 , n2800 , n2801 , n2802 , n2803 , n2805 , 
n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , 
n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2826 , n2827 , 
n2828 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , 
n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2848 , n2849 , n2850 , 
n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
n2861 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , 
n2872 , n2874 , n2875 , n2876 , n2877 , n2879 , n2880 , n2881 , n2882 , n2885 , 
n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , 
n2896 , n2897 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2926 , n2927 , n2928 , 
n2929 , n2930 , n2931 , n2932 , n2933 , n2935 , n2936 , n2937 , n2938 , n2940 , 
n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
n2961 , n2962 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , 
n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , 
n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , 
n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , 
n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , 
n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , 
n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , 
n3032 , n3033 , n3034 , n3035 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
n3043 , n3044 , n3045 , n3046 , n3047 , n3049 , n3050 , n3051 , n3052 , n3053 , 
n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , 
n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , 
n3074 , n3075 , n3077 , n3078 , n3079 , n3081 , n3082 , n3083 , n3085 , n3086 , 
n3087 , n3088 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , 
n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3107 , n3109 , n3110 , 
n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3140 , n3141 , n3142 , 
n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3164 , 
n3165 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , 
n3176 , n3177 , n3178 , n3180 , n3181 , n3182 , n3183 , n3184 , n3186 , n3187 , 
n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , 
n3198 , n3199 , n3200 , n3201 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , 
n3209 , n3210 , n3211 , n3212 , n3213 , n3215 , n3216 , n3217 , n3218 , n3219 , 
n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3229 , n3230 , 
n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , 
n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3260 , n3261 , n3262 , 
n3263 , n3264 , n3265 , n3266 , n3267 , n3269 , n3271 , n3272 , n3273 , n3274 , 
n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3283 , n3284 , n3285 , n3286 , 
n3287 , n3288 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3298 , 
n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3308 , n3309 , 
n3310 , n3311 , n3313 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , 
n3322 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , 
n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
n3343 , n3344 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , 
n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , 
n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , 
n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , 
n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3391 , n3392 , n3393 , n3395 , 
n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , 
n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , 
n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3426 , 
n3427 , n3428 , n3429 , n3430 , n3431 , n3434 , n3435 , n3436 , n3437 , n3438 , 
n3439 , n3441 , n3442 , n3443 , n3444 , n3445 , n3447 , n3448 , n3449 , n3450 , 
n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3461 , 
n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3470 , n3471 , n3472 , 
n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
n3483 , n3484 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , 
n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , 
n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , 
n3514 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3524 , n3525 , 
n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3554 , n3555 , n3556 , n3558 , 
n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , 
n3569 , n3570 , n3571 , n3572 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
n3590 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3600 , n3601 , 
n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , 
n3613 , n3615 , n3616 , n3617 , n3618 , n3619 , n3621 , n3622 , n3623 , n3625 , 
n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , 
n3636 , n3637 , n3638 , n3639 , n3640 , n3642 , n3643 , n3644 , n3645 , n3647 , 
n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , 
n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , 
n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , 
n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3687 , n3689 , 
n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3718 , n3719 , n3720 , 
n3721 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , 
n3732 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
n3753 , n3754 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , 
n3764 , n3766 , n3767 , n3768 , n3770 , n3771 , n3773 , n3774 , n3775 , n3776 , 
n3777 , n3779 , n3780 , n3781 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , 
n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , 
n3799 , n3800 , n3801 , n3802 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
n3821 , n3823 , n3824 , n3825 , n3826 , n3827 , n3829 , n3830 , n3831 , n3832 , 
n3833 , n3834 , n3835 , n3836 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , 
n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , 
n3854 , n3855 , n3856 , n3857 , n3859 , n3860 , n3861 , n3862 , n3864 , n3865 , 
n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , 
n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , 
n3886 , n3887 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3918 , 
n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3929 , 
n3930 , n3931 , n3932 , n3933 , n3934 , n3936 , n3938 , n3939 , n3940 , n3941 , 
n3943 , n3944 , n3945 , n3946 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , 
n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , 
n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , 
n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3982 , n3983 , n3984 , 
n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3997 , n3998 , 
n3999 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
n4010 , n4011 , n4012 , n4013 , n4014 , n4016 , n4017 , n4018 , n4019 , n4020 , 
n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
n4031 , n4032 , n4033 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , 
n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4052 , 
n4053 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , 
n4064 , n4065 , n4066 , n4067 , n4068 , n4070 , n4071 , n4072 , n4074 , n4075 , 
n4076 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4096 , n4097 , 
n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , 
n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , 
n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , 
n4128 , n4129 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
n4189 , n4191 , n4192 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
n4211 , n4212 , n4214 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , 
n4223 , n4224 , n4225 , n4226 , n4227 , n4229 , n4230 , n4231 , n4232 , n4233 , 
n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , 
n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , 
n4254 , n4255 , n4256 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , 
n4265 , n4266 , n4267 , n4268 , n4269 , n4271 , n4272 , n4273 , n4274 , n4275 , 
n4276 , n4277 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
n4297 , n4298 , n4299 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , 
n4308 , n4309 , n4310 , n4311 , n4312 , n4314 , n4315 , n4316 , n4318 , n4319 , 
n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
n4330 , n4331 , n4332 , n4333 , n4334 , n4336 , n4337 , n4338 , n4339 , n4340 , 
n4341 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4351 , n4352 , 
n4353 , n4354 , n4355 , n4356 , n4357 , n4359 , n4360 , n4361 , n4362 , n4363 , 
n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , 
n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , 
n4384 , n4385 , n4386 , n4387 , n4389 , n4390 , n4391 , n4392 , n4394 , n4395 , 
n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , 
n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , 
n4416 , n4417 , n4418 , n4420 , n4421 , n4423 , n4424 , n4425 , n4426 , n4427 , 
n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , 
n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , 
n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , 
n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , 
n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , 
n4478 , n4479 , n4480 , n4481 , n4483 , n4484 , n4485 , n4486 , n4488 , n4489 , 
n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
n4510 , n4511 , n4512 , n4513 , n4514 , n4516 , n4517 , n4518 , n4519 , n4520 , 
n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4531 , n4532 , 
n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , 
n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , 
n4553 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , 
n4564 , n4565 , n4566 , n4567 , n4568 , n4570 , n4571 , n4572 , n4573 , n4574 , 
n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , 
n4595 , n4596 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , 
n4606 , n4607 , n4608 , n4609 , n4610 , n4612 , n4613 , n4614 , n4615 , n4616 , 
n4617 , n4618 , n4619 , n4621 , n4623 , n4624 , n4626 , n4627 , n4628 , n4629 , 
n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
n4640 , n4641 , n4643 , n4644 , n4645 , n4646 , n4648 , n4649 , n4650 , n4651 , 
n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , 
n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , 
n4673 , n4674 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , 
n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , 
n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , 
n4704 , n4705 , n4706 , n4707 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , 
n4715 , n4716 , n4717 , n4718 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , 
n4726 , n4728 , n4729 , n4730 , n4731 , n4732 , n4734 , n4735 , n4737 , n4738 , 
n4739 , n4740 , n4741 , n4742 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
n4770 , n4771 , n4772 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
n4781 , n4782 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , 
n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , 
n4802 , n4803 , n4804 , n4806 , n4807 , n4808 , n4809 , n4811 , n4812 , n4813 , 
n4814 , n4815 , n4816 , n4817 , n4818 , n4820 , n4821 , n4822 , n4823 , n4824 , 
n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , 
n4835 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4845 , n4846 , 
n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , 
n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , 
n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , 
n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , 
n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , 
n4898 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
n4919 , n4921 , n4922 , n4923 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
n4931 , n4932 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , 
n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , 
n4952 , n4953 , n4954 , n4955 , n4957 , n4960 , n4961 , n4962 , n4963 , n4964 , 
n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , 
n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , 
n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , 
n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5004 , n5005 , 
n5006 , n5007 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
n5017 , n5018 , n5019 , n5020 , n5021 , n5023 , n5025 , n5026 , n5027 , n5028 , 
n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
n5049 , n5050 , n5051 , n5052 , n5053 , n5055 , n5056 , n5057 , n5058 , n5059 , 
n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5070 , 
n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5089 , n5090 , n5091 , 
n5092 , n5093 , n5094 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , 
n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , 
n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , 
n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , 
n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , 
n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5151 , n5152 , n5153 , n5154 , 
n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5165 , 
n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , 
n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , 
n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , 
n5196 , n5197 , n5198 , n5199 , n5200 , n5202 , n5203 , n5204 , n5205 , n5206 , 
n5207 , n5208 , n5209 , n5210 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5227 , n5228 , n5229 , 
n5230 , n5231 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
n5241 , n5242 , n5243 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5252 , 
n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , 
n5263 , n5264 , n5265 , n5266 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , 
n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , 
n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , 
n5294 , n5296 , n5297 , n5298 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5314 , n5315 , n5316 , n5317 , 
n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , 
n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , 
n5338 , n5339 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
n5372 , n5373 , n5374 , n5375 , n5376 , n5378 , n5379 , n5380 , n5381 , n5382 , 
n5383 , n5384 , n5386 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , 
n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , 
n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , 
n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , 
n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , 
n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5443 , n5444 , n5445 , n5446 , 
n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
n5477 , n5478 , n5479 , n5480 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , 
n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , 
n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , 
n5508 , n5509 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
n5580 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
n5591 , n5592 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , 
n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , 
n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , 
n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , 
n5632 , n5634 , n5635 , n5637 , n5639 , n5641 , n5642 , n5644 , n5645 , n5646 , 
n5647 , n5648 , n5650 , n5651 , n5652 , n5653 , n5654 , n5656 , n5657 , n5658 , 
n5659 , n5660 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5669 , n5671 , 
n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , 
n5682 , n5683 , n5684 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , 
n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , 
n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , 
n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5722 , n5723 , 
n5724 , n5725 , n5726 , n5728 , n5729 , n5730 , n5731 , n5733 , n5734 , n5735 , 
n5736 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
n5757 , n5758 , n5759 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , 
n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , 
n5778 , n5779 , n5780 , n5781 , n5782 , n5784 , n5785 , n5786 , n5787 , n5788 , 
n5789 , n5790 , n5791 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
n5830 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
n5871 , n5872 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , 
n5882 , n5883 , n5884 , n5885 , n5887 , n5889 , n5890 , n5891 , n5892 , n5893 , 
n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5904 , 
n5905 , n5906 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , 
n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5923 , n5924 , n5925 , n5926 , 
n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
n5938 , n5939 , n5940 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5949 , 
n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5958 , n5959 , n5960 , 
n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
n6031 , n6032 , n6033 , n6034 , n6035 , n6037 , n6038 , n6040 , n6041 , n6042 , 
n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , 
n6053 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , 
n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , 
n6075 , n6076 , n6077 , n6078 , n6079 , n6081 , n6082 , n6083 , n6084 , n6085 , 
n6086 , n6087 , n6088 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6106 , n6107 , 
n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6115 , n6116 , n6117 , n6118 , 
n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6128 , n6129 , 
n6130 , n6131 , n6132 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
n6142 , n6143 , n6144 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , 
n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , 
n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6173 , 
n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , 
n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , 
n6195 , n6197 , n6198 , n6199 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , 
n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , 
n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6224 , n6225 , n6226 , n6227 , 
n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , 
n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , 
n6248 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6257 , n6258 , n6260 , 
n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
n6291 , n6292 , n6293 , n6294 , n6296 , n6297 , n6299 , n6300 , n6301 , n6302 , 
n6303 , n6304 , n6305 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6314 , 
n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , 
n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6332 , n6333 , n6335 , n6336 , 
n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , 
n6348 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
n6359 , n6360 , n6361 , n6363 , n6364 , n6365 , n6367 , n6368 , n6369 , n6370 , 
n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6391 , 
n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , 
n6402 , n6404 , n6405 , n6406 , n6407 , n6408 , n6410 , n6411 , n6412 , n6413 , 
n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , 
n6424 , n6425 , n6426 , n6428 , n6429 , n6432 , n6433 , n6434 , n6435 , n6436 , 
n6437 , n6438 , n6439 , n6441 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
n6449 , n6450 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6459 , n6460 , 
n6461 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6471 , n6472 , 
n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , 
n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , 
n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , 
n6503 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , 
n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , 
n6525 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6535 , n6536 , n6537 , 
n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6545 , n6547 , n6548 , n6549 , 
n6550 , n6551 , n6552 , n6553 , n6554 , n6556 , n6557 , n6558 , n6559 , n6560 , 
n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
n6601 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , 
n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , 
n6623 , n6624 , n6625 , n6627 , n6628 , n6629 , n6630 , n6631 , n6633 , n6634 , 
n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6652 , n6653 , n6654 , n6655 , 
n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , 
n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , 
n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , 
n6686 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
n6707 , n6708 , n6709 , n6710 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , 
n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , 
n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6735 , n6736 , n6737 , n6738 , 
n6739 , n6740 , n6741 , n6742 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
n6790 , n6791 , n6792 , n6793 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
n6801 , n6802 , n6804 , n6805 , n6806 , n6807 , n6808 , n6810 , n6811 , n6812 , 
n6814 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6863 , n6864 , n6865 , 
n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6875 , n6876 , 
n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
n6887 , n6889 , n6890 , n6891 , n6892 , n6894 , n6895 , n6896 , n6897 , n6898 , 
n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
n6941 , n6942 , n6943 , n6944 , n6945 , n6947 , n6948 , n6949 , n6950 , n6951 , 
n6952 , n6953 , n6954 , n6955 , n6956 , n6958 , n6959 , n6960 , n6961 , n6962 , 
n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , 
n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
n6983 , n6984 , n6985 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , 
n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , 
n7004 , n7005 , n7006 , n7007 , n7008 , n7010 , n7011 , n7012 , n7013 , n7015 , 
n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7025 , n7026 , n7027 , 
n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , 
n7038 , n7039 , n7040 , n7041 , n7042 , n7044 , n7045 , n7048 , n7049 , n7050 , 
n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
n7071 , n7072 , n7073 , n7074 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , 
n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , 
n7093 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , 
n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , 
n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , 
n7124 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
n7145 , n7146 , n7147 , n7149 , n7151 , n7152 , n7153 , n7154 , n7156 , n7157 , 
n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , 
n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , 
n7178 , n7179 , n7181 , n7182 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7211 , n7212 , 
n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , 
n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7232 , n7233 , 
n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7242 , n7243 , n7244 , 
n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7266 , 
n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , 
n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , 
n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
n7309 , n7310 , n7311 , n7312 , n7313 , n7316 , n7317 , n7318 , n7319 , n7320 , 
n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
n7341 , n7342 , n7343 , n7344 , n7345 , n7347 , n7348 , n7349 , n7350 , n7351 , 
n7352 , n7353 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , 
n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7372 , n7373 , n7374 , 
n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
n7385 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , 
n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , 
n7406 , n7407 , n7408 , n7409 , n7410 , n7412 , n7413 , n7415 , n7416 , n7417 , 
n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7426 , n7427 , n7429 , 
n7430 , n7431 , n7432 , n7433 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7448 , n7449 , n7450 , n7451 , 
n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , 
n7462 , n7463 , n7464 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , 
n7474 , n7475 , n7476 , n7477 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , 
n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7503 , n7504 , n7505 , n7506 , 
n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
n7537 , n7538 , n7539 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , 
n7548 , n7549 , n7550 , n7551 , n7552 , n7554 , n7555 , n7556 , n7557 , n7558 , 
n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
n7589 , n7590 , n7591 , n7592 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
n7650 , n7652 , n7653 , n7654 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , 
n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7669 , n7670 , n7671 , n7672 , 
n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , 
n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7693 , 
n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7702 , n7703 , n7704 , 
n7706 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , 
n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , 
n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7736 , n7737 , n7738 , n7739 , 
n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , 
n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , 
n7782 , n7783 , n7784 , n7785 , n7786 , n7788 , n7789 , n7790 , n7791 , n7792 , 
n7793 , n7794 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , 
n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , 
n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , 
n7824 , n7825 , n7826 , n7827 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7853 , n7854 , n7855 , 
n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7863 , n7864 , n7865 , n7866 , 
n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
n7877 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , 
n7888 , n7889 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7949 , 
n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7988 , n7989 , n7990 , 
n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
n8001 , n8002 , n8003 , n8004 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , 
n8012 , n8013 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , 
n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8031 , n8032 , n8033 , 
n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8043 , n8044 , 
n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8064 , n8065 , 
n8066 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8077 , 
n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , 
n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8096 , n8098 , n8099 , 
n8100 , n8101 , n8102 , n8103 , n8105 , n8106 , n8107 , n8108 , n8110 , n8111 , 
n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , 
n8122 , n8123 , n8124 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , 
n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , 
n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , 
n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , 
n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , 
n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8181 , n8182 , n8184 , 
n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8195 , 
n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , 
n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , 
n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , 
n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8236 , 
n8237 , n8238 , n8239 , n8240 , n8241 , n8243 , n8244 , n8245 , n8246 , n8247 , 
n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , 
n8258 , n8259 , n8261 , n8262 , n8263 , n8265 , n8266 , n8267 , n8268 , n8269 , 
n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
n8291 , n8292 , n8293 , n8294 , n8295 , n8298 , n8299 , n8300 , n8302 , n8303 , 
n8304 , n8305 , n8306 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8315 , 
n8316 , n8317 , n8318 , n8322 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
n8360 , n8361 , n8362 , n8363 , n8364 , n8366 , n8367 , n8368 , n8369 , n8370 , 
n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8381 , n8382 , 
n8383 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , 
n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , 
n8404 , n8405 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , 
n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , 
n8426 , n8427 , n8428 , n8429 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
n8457 , n8458 , n8459 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , 
n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , 
n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8486 , n8487 , n8488 , 
n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
n8509 , n8510 , n8511 , n8512 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
n8560 , n8562 , n8563 , n8564 , n8565 , n8567 , n8568 , n8569 , n8571 , n8572 , 
n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , 
n8583 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , 
n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , 
n8604 , n8605 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , 
n8615 , n8616 , n8617 , n8618 , n8619 , n8622 , n8623 , n8624 , n8625 , n8626 , 
n8627 , n8629 , n8630 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8686 , n8687 , n8688 , n8690 , 
n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
n8701 , n8702 , n8703 , n8704 , n8705 , n8707 , n8708 , n8709 , n8710 , n8711 , 
n8712 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , 
n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , 
n8734 , n8735 , n8736 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , 
n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , 
n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , 
n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8772 , n8773 , n8774 , n8775 , 
n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8785 , n8786 , 
n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8805 , n8806 , n8807 , 
n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
n8819 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
n8830 , n8831 , n8832 , n8833 , n8835 , n8837 , n8838 , n8839 , n8840 , n8841 , 
n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , 
n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , 
n8862 , n8863 , n8864 , n8865 , n8866 , n8868 , n8869 , n8870 , n8871 , n8872 , 
n8874 , n8875 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , 
n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , 
n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8903 , n8904 , n8905 , 
n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , 
n8916 , n8917 , n8918 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
n8947 , n8948 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , 
n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8987 , n8989 , n8990 , 
n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , 
n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , 
n9032 , n9033 , n9034 , n9035 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , 
n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , 
n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , 
n9064 , n9065 , n9066 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , 
n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , 
n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , 
n9095 , n9096 , n9097 , n9098 , n9100 , n9101 , n9102 , n9103 , n9104 , n9106 , 
n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9117 , n9118 , 
n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
n9129 , n9130 , n9131 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
n9140 , n9141 , n9142 , n9143 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , 
n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , 
n9162 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , 
n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , 
n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , 
n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , 
n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9210 , n9211 , n9212 , n9213 , 
n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9224 , 
n9225 , n9226 , n9227 , n9229 , n9230 , n9231 , n9232 , n9233 , n9235 , n9236 , 
n9237 , n9238 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9247 , n9248 , 
n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9259 , 
n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
n9270 , n9271 , n9272 , n9273 , n9275 , n9276 , n9278 , n9279 , n9280 , n9281 , 
n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , 
n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , 
n9302 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9311 , n9312 , n9313 , 
n9314 , n9315 , n9316 , n9317 , n9319 , n9320 , n9322 , n9323 , n9324 , n9325 , 
n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , 
n9337 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , 
n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , 
n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
n9409 , n9410 , n9411 , n9412 , n9413 , n9415 , n9416 , n9417 , n9418 , n9419 , 
n9420 , n9421 , n9422 , n9423 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9470 , n9471 , 
n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , 
n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , 
n9492 , n9493 , n9494 , n9495 , n9496 , n9498 , n9499 , n9500 , n9501 , n9502 , 
n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9510 , n9511 , n9512 , n9513 , 
n9514 , n9515 , n9516 , n9518 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , 
n9527 , n9528 , n9529 , n9530 , n9531 , n9533 , n9534 , n9536 , n9537 , n9538 , 
n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
n9549 , n9550 , n9551 , n9552 , n9553 , n9555 , n9556 , n9557 , n9558 , n9559 , 
n9560 , n9561 , n9562 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
n9592 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , 
n9603 , n9605 , n9606 , n9607 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
n9615 , n9616 , n9617 , n9618 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , 
n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9633 , n9634 , n9635 , n9636 , 
n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9644 , n9645 , n9646 , n9648 , 
n9649 , n9650 , n9651 , n9652 , n9654 , n9657 , n9658 , n9659 , n9660 , n9661 , 
n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , 
n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , 
n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9692 , 
n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , 
n9703 , n9704 , n9705 , n9706 , n9707 , n9709 , n9710 , n9711 , n9712 , n9713 , 
n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , 
n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , 
n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , 
n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , 
n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , 
n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , 
n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , 
n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , 
n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
n9827 , n9828 , n9829 , n9830 , n9832 , n9833 , n9834 , n9836 , n9837 , n9838 , 
n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
n9849 , n9850 , n9851 , n9852 , n9853 , n9855 , n9856 , n9857 , n9858 , n9859 , 
n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9899 , n9900 , n9901 , 
n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9909 , n9910 , n9911 , n9912 , 
n9913 , n9914 , n9915 , n9916 , n9917 , n9919 , n9920 , n9921 , n9922 , n9923 , 
n9924 , n9925 , n9926 , n9927 , n9928 , n9930 , n9931 , n9932 , n9933 , n9934 , 
n9936 , n9937 , n9938 , n9940 , n9941 , n9942 , n9943 , n9944 , n9946 , n9947 , 
n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
n9981 , n9982 , n9983 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , 
n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , 
n10003 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , 
n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , 
n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10035 , 
n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , 
n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , 
n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , 
n10066 , n10067 , n10068 , n10069 , n10070 , n10072 , n10073 , n10074 , n10075 , n10076 , 
n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , 
n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10096 , n10097 , n10098 , 
n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
n10109 , n10110 , n10111 , n10112 , n10113 , n10115 , n10116 , n10118 , n10119 , n10120 , 
n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10129 , n10130 , n10131 , n10132 , 
n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10141 , n10142 , n10143 , n10144 , 
n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , 
n10155 , n10157 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
n10167 , n10168 , n10169 , n10170 , n10173 , n10175 , n10177 , n10178 , n10179 , n10180 , 
n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
n10191 , n10192 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , 
n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10210 , n10211 , n10212 , 
n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , 
n10223 , n10224 , n10225 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , 
n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , 
n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10252 , n10253 , n10255 , 
n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10264 , n10265 , n10266 , 
n10267 , n10268 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , 
n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , 
n10288 , n10289 , n10290 , n10291 , n10293 , n10294 , n10295 , n10297 , n10298 , n10299 , 
n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10307 , n10308 , n10309 , n10310 , 
n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10321 , 
n10322 , n10323 , n10324 , n10325 , n10326 , n10328 , n10329 , n10330 , n10331 , n10332 , 
n10333 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , 
n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10354 , n10355 , n10356 , 
n10357 , n10359 , n10360 , n10361 , n10362 , n10364 , n10366 , n10367 , n10368 , n10369 , 
n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
n10390 , n10391 , n10392 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , 
n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10409 , n10410 , n10411 , 
n10412 , n10414 , n10415 , n10416 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , 
n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10434 , 
n10435 , n10436 , n10437 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , 
n10446 , n10447 , n10448 , n10449 , n10450 , n10452 , n10453 , n10454 , n10455 , n10456 , 
n10457 , n10458 , n10459 , n10460 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , 
n10468 , n10469 , n10470 , n10472 , n10473 , n10476 , n10478 , n10479 , n10480 , n10481 , 
n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10491 , n10492 , 
n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , 
n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , 
n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10522 , n10523 , 
n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , 
n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , 
n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10552 , n10554 , n10555 , 
n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , 
n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , 
n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10584 , n10585 , n10586 , 
n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10616 , n10617 , 
n10618 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
n10641 , n10642 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , 
n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , 
n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , 
n10672 , n10673 , n10674 , n10675 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , 
n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10691 , n10693 , n10694 , 
n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , 
n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , 
n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , 
n10725 , n10726 , n10727 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , 
n10736 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10754 , n10755 , n10756 , n10757 , 
n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , 
n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , 
n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , 
n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10796 , n10797 , n10798 , 
n10799 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
n10820 , n10821 , n10822 , n10823 , n10824 , n10826 , n10827 , n10828 , n10829 , n10830 , 
n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , 
n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , 
n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , 
n10861 , n10862 , n10863 , n10864 , n10867 , n10869 , n10870 , n10871 , n10872 , n10873 , 
n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , 
n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , 
n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , 
n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10911 , n10912 , n10913 , n10915 , 
n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , 
n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , 
n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , 
n10946 , n10947 , n10948 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10957 , 
n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10967 , n10968 , 
n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10978 , n10979 , 
n10980 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10991 , 
n10992 , n10993 , n10994 , n10995 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , 
n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , 
n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , 
n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11032 , n11033 , n11034 , 
n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , 
n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11052 , n11053 , n11054 , n11055 , 
n11056 , n11057 , n11058 , n11059 , n11061 , n11063 , n11064 , n11066 , n11067 , n11068 , 
n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
n11129 , n11130 , n11131 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , 
n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , 
n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , 
n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , 
n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , 
n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11198 , n11199 , n11200 , n11201 , 
n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11209 , n11210 , n11211 , n11212 , 
n11213 , n11214 , n11215 , n11216 , n11217 , n11219 , n11220 , n11221 , n11222 , n11224 , 
n11225 , n11226 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , 
n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11246 , 
n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11254 , n11255 , n11256 , n11257 , 
n11258 , n11259 , n11260 , n11261 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11329 , n11330 , 
n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11339 , n11340 , n11341 , 
n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , 
n11352 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11362 , n11363 , n11364 , 
n11365 , n11366 , n11367 , n11369 , n11370 , n11371 , n11372 , n11374 , n11375 , n11376 , 
n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
n11397 , n11398 , n11399 , n11400 , n11402 , n11403 , n11404 , n11405 , n11406 , n11408 , 
n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
n11429 , n11430 , n11431 , n11432 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
n11460 , n11461 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , 
n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , 
n11481 , n11482 , n11483 , n11484 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , 
n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , 
n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , 
n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , 
n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , 
n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , 
n11542 , n11543 , n11544 , n11545 , n11546 , n11548 , n11549 , n11550 , n11551 , n11552 , 
n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , 
n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , 
n11573 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , 
n11584 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , 
n11595 , n11596 , n11597 , n11598 , n11600 , n11602 , n11603 , n11604 , n11605 , n11606 , 
n11607 , n11608 , n11609 , n11611 , n11612 , n11615 , n11616 , n11617 , n11618 , n11619 , 
n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
n11630 , n11631 , n11632 , n11633 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , 
n11641 , n11642 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , 
n11652 , n11654 , n11655 , n11656 , n11657 , n11659 , n11660 , n11661 , n11662 , n11663 , 
n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , 
n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11683 , n11684 , 
n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11693 , n11694 , n11695 , n11696 , 
n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
n11707 , n11708 , n11709 , n11710 , n11712 , n11713 , n11715 , n11716 , n11717 , n11718 , 
n11719 , n11720 , n11721 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11737 , n11738 , n11739 , n11740 , 
n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , 
n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , 
n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , 
n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , 
n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11790 , n11791 , n11793 , 
n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , 
n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11813 , n11815 , 
n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , 
n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , 
n11836 , n11837 , n11838 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11848 , 
n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11867 , n11868 , n11869 , 
n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
n11880 , n11881 , n11882 , n11883 , n11885 , n11887 , n11888 , n11889 , n11890 , n11891 , 
n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , 
n11902 , n11903 , n11904 , n11906 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , 
n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , 
n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , 
n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , 
n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , 
n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11964 , 
n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , 
n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11985 , 
n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , 
n11996 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12025 , n12026 , n12027 , 
n12028 , n12029 , n12031 , n12033 , n12034 , n12036 , n12037 , n12039 , n12040 , n12041 , 
n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12050 , n12051 , n12052 , 
n12053 , n12054 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , 
n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12073 , n12074 , 
n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , 
n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , 
n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , 
n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , 
n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , 
n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12136 , n12137 , n12138 , 
n12139 , n12140 , n12141 , n12142 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
n12160 , n12161 , n12162 , n12163 , n12164 , n12166 , n12167 , n12168 , n12169 , n12170 , 
n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , 
n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , 
n12192 , n12193 , n12195 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , 
n12204 , n12205 , n12206 , n12208 , n12209 , n12211 , n12212 , n12213 , n12214 , n12215 , 
n12216 , n12217 , n12218 , n12219 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
n12227 , n12228 , n12229 , n12230 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , 
n12238 , n12239 , n12240 , n12241 , n12244 , n12246 , n12247 , n12248 , n12249 , n12250 , 
n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12260 , n12261 , 
n12262 , n12263 , n12264 , n12266 , n12267 , n12268 , n12269 , n12270 , n12272 , n12273 , 
n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , 
n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , 
n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , 
n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12313 , n12314 , 
n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , 
n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , 
n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , 
n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , 
n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12365 , 
n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12375 , n12376 , 
n12377 , n12378 , n12379 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , 
n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , 
n12400 , n12401 , n12402 , n12403 , n12405 , n12406 , n12407 , n12408 , n12410 , n12411 , 
n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , 
n12422 , n12423 , n12424 , n12425 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , 
n12433 , n12434 , n12435 , n12436 , n12437 , n12439 , n12440 , n12441 , n12442 , n12443 , 
n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , 
n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12465 , 
n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , 
n12476 , n12477 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12496 , n12497 , 
n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , 
n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12515 , n12516 , n12517 , n12518 , 
n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , 
n12529 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
n12560 , n12562 , n12563 , n12564 , n12565 , n12567 , n12568 , n12569 , n12570 , n12571 , 
n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , 
n12583 , n12584 , n12585 , n12586 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , 
n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , 
n12604 , n12606 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , 
n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12626 , 
n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , 
n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , 
n12649 , n12650 , n12651 , n12652 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12670 , n12671 , 
n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12679 , n12680 , n12682 , n12683 , 
n12684 , n12685 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , 
n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12705 , n12706 , 
n12708 , n12709 , n12710 , n12711 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12727 , n12728 , n12729 , n12730 , 
n12731 , n12732 , n12733 , n12735 , n12736 , n12738 , n12739 , n12740 , n12741 , n12742 , 
n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , 
n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , 
n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , 
n12773 , n12774 , n12775 , n12776 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , 
n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , 
n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12804 , 
n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12815 , n12816 , n12817 , 
n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , 
n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , 
n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , 
n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , 
n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , 
n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , 
n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12921 , 
n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , 
n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , 
n12943 , n12944 , n12945 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , 
n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , 
n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , 
n12974 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , 
n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , 
n12995 , n12996 , n12997 , n12999 , n13000 , n13001 , n13002 , n13003 , n13005 , n13006 , 
n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
n13017 , n13018 , n13019 , n13020 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , 
n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , 
n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , 
n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
n13059 , n13060 , n13061 , n13062 , n13063 , n13065 , n13066 , n13067 , n13068 , n13069 , 
n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
n13100 , n13101 , n13102 , n13103 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , 
n13111 , n13112 , n13113 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , 
n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , 
n13132 , n13133 , n13134 , n13135 , n13136 , n13138 , n13139 , n13140 , n13141 , n13142 , 
n13143 , n13144 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , 
n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13162 , n13163 , n13164 , 
n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , 
n13175 , n13176 , n13177 , n13178 , n13180 , n13182 , n13183 , n13184 , n13185 , n13186 , 
n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
n13207 , n13208 , n13209 , n13212 , n13213 , n13214 , n13216 , n13217 , n13218 , n13220 , 
n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , 
n13231 , n13232 , n13233 , n13236 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , 
n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , 
n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , 
n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13272 , n13273 , n13274 , 
n13275 , n13277 , n13278 , n13279 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
n13287 , n13288 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , 
n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , 
n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , 
n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , 
n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , 
n13339 , n13340 , n13341 , n13342 , n13343 , n13346 , n13347 , n13348 , n13349 , n13350 , 
n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13359 , n13361 , n13362 , 
n13363 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13375 , 
n13376 , n13377 , n13378 , n13379 , n13381 , n13382 , n13383 , n13384 , n13386 , n13387 , 
n13388 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , 
n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13407 , n13408 , n13409 , n13411 , 
n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , 
n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , 
n13432 , n13433 , n13434 , n13435 , n13436 , n13438 , n13439 , n13440 , n13441 , n13442 , 
n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13451 , n13452 , n13455 , 
n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , 
n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , 
n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , 
n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13495 , n13496 , 
n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13505 , n13506 , n13507 , 
n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13515 , n13516 , n13517 , n13518 , 
n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13527 , n13528 , n13529 , 
n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
n13540 , n13541 , n13542 , n13543 , n13544 , n13546 , n13547 , n13548 , n13549 , n13550 , 
n13551 , n13552 , n13553 , n13554 , n13555 , n13557 , n13558 , n13560 , n13561 , n13563 , 
n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , 
n13574 , n13575 , n13576 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , 
n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , 
n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13605 , 
n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , 
n13616 , n13617 , n13618 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13636 , n13637 , 
n13638 , n13639 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
n13649 , n13650 , n13651 , n13652 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , 
n13662 , n13663 , n13664 , n13665 , n13666 , n13668 , n13669 , n13670 , n13671 , n13672 , 
n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13680 , n13681 , n13682 , n13683 , 
n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , 
n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13702 , n13703 , n13704 , n13705 , 
n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , 
n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13726 , 
n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
n13747 , n13748 , n13749 , n13750 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , 
n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , 
n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , 
n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , 
n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , 
n13798 , n13799 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13809 , 
n13810 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , 
n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , 
n13831 , n13832 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , 
n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13851 , n13852 , n13853 , 
n13854 , n13855 , n13856 , n13857 , n13858 , n13860 , n13862 , n13863 , n13864 , n13865 , 
n13866 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
n13907 , n13908 , n13909 , n13911 , n13912 , n13913 , n13915 , n13916 , n13917 , n13918 , 
n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , 
n13929 , n13930 , n13931 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , 
n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , 
n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13958 , n13959 , n13960 , 
n13961 , n13962 , n13963 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , 
n13972 , n13973 , n13974 , n13976 , n13977 , n13978 , n13979 , n13981 , n13982 , n13983 , 
n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , 
n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , 
n14005 , n14006 , n14007 , n14009 , n14010 , n14011 , n14013 , n14014 , n14015 , n14017 , 
n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , 
n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14036 , n14037 , n14038 , n14039 , 
n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14050 , n14051 , 
n14052 , n14053 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , 
n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , 
n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , 
n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , 
n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , 
n14104 , n14105 , n14107 , n14108 , n14109 , n14111 , n14113 , n14114 , n14115 , n14116 , 
n14117 , n14118 , n14119 , n14120 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , 
n14128 , n14129 , n14130 , n14132 , n14133 , n14134 , n14135 , n14138 , n14139 , n14140 , 
n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , 
n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , 
n14161 , n14162 , n14163 , n14164 , n14165 , n14168 , n14169 , n14170 , n14171 , n14172 , 
n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , 
n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , 
n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14201 , n14202 , n14203 , 
n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14213 , n14214 , 
n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , 
n14225 , n14226 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , 
n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , 
n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , 
n14256 , n14257 , n14258 , n14260 , n14261 , n14263 , n14264 , n14265 , n14266 , n14267 , 
n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , 
n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , 
n14288 , n14289 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , 
n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , 
n14309 , n14310 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , 
n14320 , n14321 , n14322 , n14323 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , 
n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , 
n14341 , n14342 , n14343 , n14345 , n14346 , n14347 , n14349 , n14350 , n14351 , n14352 , 
n14353 , n14354 , n14355 , n14357 , n14358 , n14359 , n14360 , n14362 , n14364 , n14365 , 
n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , 
n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , 
n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , 
n14396 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
n14407 , n14408 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , 
n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , 
n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14436 , n14437 , n14438 , n14439 , 
n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , 
n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14478 , n14479 , n14480 , 
n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14491 , n14492 , 
n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , 
n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , 
n14515 , n14516 , n14517 , n14518 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
n14527 , n14528 , n14529 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , 
n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , 
n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14556 , n14557 , n14558 , 
n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14566 , n14567 , n14568 , n14569 , 
n14570 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , 
n14581 , n14582 , n14583 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , 
n14592 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , 
n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14614 , 
n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14625 , 
n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , 
n14636 , n14637 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14656 , n14657 , 
n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14666 , n14667 , n14668 , 
n14669 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , 
n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , 
n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14700 , n14701 , 
n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14712 , 
n14713 , n14714 , n14715 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , 
n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , 
n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , 
n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14754 , 
n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , 
n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , 
n14775 , n14776 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , 
n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14793 , n14794 , n14796 , n14797 , 
n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , 
n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , 
n14818 , n14819 , n14820 , n14821 , n14823 , n14824 , n14825 , n14827 , n14829 , n14830 , 
n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14838 , n14839 , n14840 , n14841 , 
n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , 
n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , 
n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , 
n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14881 , n14882 , n14884 , 
n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
n14905 , n14906 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , 
n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14926 , 
n14927 , n14929 , n14930 , n14931 , n14932 , n14933 , n14935 , n14936 , n14937 , n14938 , 
n14939 , n14940 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , 
n14950 , n14951 , n14952 , n14953 , n14955 , n14956 , n14957 , n14959 , n14960 , n14961 , 
n14963 , n14964 , n14965 , n14966 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , 
n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , 
n14984 , n14986 , n14987 , n14988 , n14990 , n14991 , n14993 , n14994 , n14995 , n14996 , 
n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
n15008 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , 
n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15027 , n15028 , n15029 , n15030 , 
n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , 
n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15050 , n15051 , 
n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15060 , n15061 , n15062 , 
n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , 
n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , 
n15083 , n15084 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , 
n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15101 , n15102 , n15103 , n15104 , 
n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , 
n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , 
n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15134 , n15135 , n15136 , 
n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15144 , n15145 , n15146 , n15147 , 
n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15156 , n15157 , n15158 , n15159 , 
n15160 , n15161 , n15162 , n15163 , n15166 , n15168 , n15169 , n15170 , n15171 , n15172 , 
n15173 , n15174 , n15175 , n15176 , n15177 , n15179 , n15180 , n15181 , n15182 , n15183 , 
n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15192 , n15193 , n15194 , 
n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , 
n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , 
n15215 , n15216 , n15217 , n15218 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , 
n15226 , n15227 , n15228 , n15229 , n15230 , n15232 , n15233 , n15234 , n15235 , n15236 , 
n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , 
n15268 , n15269 , n15270 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15279 , 
n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , 
n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , 
n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , 
n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15319 , n15320 , 
n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , 
n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15339 , n15340 , n15341 , 
n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15352 , n15353 , 
n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15364 , 
n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , 
n15375 , n15376 , n15377 , n15378 , n15380 , n15381 , n15383 , n15384 , n15385 , n15386 , 
n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15397 , 
n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15407 , n15408 , 
n15410 , n15411 , n15412 , n15414 , n15415 , n15417 , n15418 , n15419 , n15420 , n15421 , 
n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , 
n15432 , n15433 , n15435 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , 
n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , 
n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , 
n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15472 , n15473 , n15474 , 
n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15485 , 
n15486 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15495 , n15496 , n15497 , 
n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15506 , n15507 , n15508 , 
n15509 , n15510 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , 
n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , 
n15530 , n15531 , n15532 , n15533 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , 
n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , 
n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15559 , n15560 , n15561 , n15562 , 
n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , 
n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15581 , n15582 , n15583 , 
n15584 , n15585 , n15586 , n15587 , n15589 , n15590 , n15593 , n15594 , n15595 , n15596 , 
n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , 
n15607 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15619 , n15620 , 
n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , 
n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , 
n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15651 , 
n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15659 , n15660 , n15661 , n15662 , 
n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , 
n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , 
n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , 
n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , 
n15745 , n15746 , n15747 , n15748 , n15750 , n15751 , n15752 , n15754 , n15755 , n15756 , 
n15757 , n15759 , n15760 , n15761 , n15762 , n15764 , n15765 , n15766 , n15767 , n15768 , 
n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , 
n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15788 , n15789 , 
n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , 
n15801 , n15802 , n15803 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , 
n15812 , n15813 , n15814 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , 
n15823 , n15824 , n15825 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , 
n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , 
n15844 , n15845 , n15846 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , 
n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , 
n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , 
n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
n15897 , n15898 , n15899 , n15901 , n15902 , n15903 , n15905 , n15906 , n15907 , n15908 , 
n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , 
n15919 , n15920 , n15921 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , 
n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15938 , n15939 , n15940 , 
n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15948 , n15949 , n15950 , n15952 , 
n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , 
n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , 
n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , 
n15983 , n15984 , n15985 , n15989 , n15990 , n15991 , n15992 , n15994 , n15996 , n15997 , 
n15998 , n16000 , n16001 , n16002 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , 
n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16020 , 
n16021 , n16022 , n16023 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , 
n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16041 , n16042 , 
n16043 , n16044 , n16045 , n16046 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , 
n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , 
n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16071 , n16072 , n16073 , n16074 , 
n16076 , n16077 , n16078 , n16079 , n16080 , n16082 , n16083 , n16084 , n16085 , n16086 , 
n16087 , n16088 , n16089 , n16090 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , 
n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16105 , n16106 , n16107 , n16108 , 
n16109 , n16110 , n16111 , n16112 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , 
n16120 , n16121 , n16122 , n16123 , n16124 , n16126 , n16127 , n16128 , n16129 , n16130 , 
n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , 
n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , 
n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , 
n16163 , n16165 , n16166 , n16167 , n16168 , n16169 , n16171 , n16172 , n16173 , n16174 , 
n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , 
n16185 , n16186 , n16188 , n16189 , n16190 , n16191 , n16193 , n16194 , n16195 , n16196 , 
n16197 , n16198 , n16199 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , 
n16208 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , 
n16219 , n16221 , n16222 , n16224 , n16225 , n16226 , n16227 , n16229 , n16230 , n16231 , 
n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16240 , n16241 , n16242 , n16243 , 
n16244 , n16245 , n16246 , n16247 , n16248 , n16250 , n16251 , n16253 , n16254 , n16255 , 
n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , 
n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16276 , 
n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16284 , n16286 , n16287 , n16288 , 
n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , 
n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16307 , n16309 , n16310 , 
n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , 
n16321 , n16322 , n16323 , n16325 , n16326 , n16327 , n16330 , n16331 , n16332 , n16333 , 
n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , 
n16345 , n16346 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , 
n16356 , n16357 , n16358 , n16359 , n16360 , n16362 , n16363 , n16364 , n16365 , n16366 , 
n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , 
n16377 , n16378 , n16379 , n16380 , n16381 , n16383 , n16384 , n16385 , n16386 , n16387 , 
n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , 
n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16407 , n16408 , 
n16409 , n16410 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , 
n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16428 , n16429 , n16430 , 
n16431 , n16432 , n16433 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16443 , 
n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , 
n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , 
n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , 
n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , 
n16484 , n16485 , n16486 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , 
n16495 , n16496 , n16497 , n16498 , n16499 , n16501 , n16502 , n16503 , n16504 , n16505 , 
n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , 
n16517 , n16518 , n16519 , n16520 , n16521 , n16523 , n16524 , n16525 , n16526 , n16527 , 
n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , 
n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , 
n16548 , n16549 , n16550 , n16551 , n16553 , n16554 , n16555 , n16556 , n16557 , n16559 , 
n16560 , n16561 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16571 , 
n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , 
n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16592 , 
n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16602 , n16603 , 
n16604 , n16605 , n16606 , n16607 , n16608 , n16610 , n16611 , n16612 , n16613 , n16614 , 
n16615 , n16616 , n16617 , n16618 , n16620 , n16621 , n16622 , n16624 , n16625 , n16626 , 
n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , 
n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , 
n16647 , n16648 , n16649 , n16650 , n16651 , n16653 , n16654 , n16655 , n16657 , n16658 , 
n16659 , n16660 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , 
n16670 , n16672 , n16673 , n16674 , n16675 , n16677 , n16678 , n16679 , n16681 , n16682 , 
n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , 
n16693 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16704 , 
n16706 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , 
n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , 
n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16738 , n16739 , 
n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , 
n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , 
n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , 
n16770 , n16771 , n16772 , n16773 , n16774 , n16776 , n16777 , n16778 , n16779 , n16780 , 
n16781 , n16782 , n16783 , n16784 , n16786 , n16787 , n16788 , n16790 , n16791 , n16792 , 
n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16800 , n16801 , n16802 , n16804 , 
n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
n16816 , n16817 , n16818 , n16819 , n16820 , n16822 , n16823 , n16825 , n16827 , n16828 , 
n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16838 , n16839 , 
n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , 
n16850 , n16851 , n16854 , n16855 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , 
n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , 
n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , 
n16884 , n16885 , n16886 , n16887 , n16889 , n16890 , n16891 , n16892 , n16894 , n16895 , 
n16896 , n16897 , n16898 , n16899 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , 
n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16917 , 
n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16928 , 
n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16938 , n16939 , 
n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , 
n16950 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
n16981 , n16982 , n16983 , n16984 , n16985 , n16987 , n16988 , n16989 , n16990 , n16991 , 
n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16999 , n17000 , n17001 , n17002 , 
n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , 
n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17020 , n17021 , n17022 , n17023 , 
n17024 , n17025 , n17026 , n17027 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , 
n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , 
n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17053 , n17054 , n17056 , n17057 , 
n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17069 , 
n17070 , n17071 , n17072 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , 
n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17090 , n17091 , 
n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , 
n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17110 , n17111 , n17112 , 
n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , 
n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , 
n17133 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , 
n17144 , n17145 , n17146 , n17147 , n17148 , n17150 , n17151 , n17152 , n17153 , n17154 , 
n17155 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , 
n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , 
n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , 
n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , 
n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , 
n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17216 , 
n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , 
n17228 , n17229 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , 
n17239 , n17240 , n17241 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , 
n17250 , n17251 , n17252 , n17253 , n17254 , n17256 , n17257 , n17258 , n17259 , n17260 , 
n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , 
n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , 
n17281 , n17282 , n17283 , n17284 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , 
n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , 
n17303 , n17304 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , 
n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , 
n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , 
n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , 
n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17355 , 
n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , 
n17366 , n17367 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , 
n17377 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , 
n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17397 , n17398 , n17399 , 
n17400 , n17401 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , 
n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17418 , n17420 , n17421 , n17422 , 
n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , 
n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17440 , n17441 , n17442 , n17443 , 
n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , 
n17455 , n17456 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , 
n17466 , n17467 , n17468 , n17469 , n17472 , n17474 , n17475 , n17476 , n17477 , n17478 , 
n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , 
n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17496 , n17497 , n17500 , n17501 , 
n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17511 , n17512 , n17513 , 
n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , 
n17525 , n17526 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , 
n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , 
n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , 
n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , 
n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , 
n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17587 , 
n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , 
n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17608 , n17609 , 
n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17618 , n17619 , n17620 , 
n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17631 , 
n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , 
n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , 
n17652 , n17653 , n17654 , n17655 , n17656 , n17658 , n17659 , n17660 , n17661 , n17662 , 
n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , 
n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , 
n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , 
n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , 
n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17713 , n17714 , n17715 , n17716 , 
n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , 
n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , 
n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17746 , n17747 , 
n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , 
n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , 
n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , 
n17779 , n17780 , n17781 , n17782 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , 
n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17799 , n17800 , 
n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17809 , n17810 , n17811 , 
n17812 , n17813 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , 
n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17830 , n17831 , n17832 , n17833 , 
n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17844 , 
n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17852 , n17853 , n17854 , n17856 , 
n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , 
n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , 
n17878 , n17879 , n17880 , n17881 , n17882 , n17884 , n17885 , n17886 , n17887 , n17888 , 
n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , 
n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , 
n17909 , n17911 , n17912 , n17913 , n17915 , n17917 , n17918 , n17919 , n17920 , n17921 , 
n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , 
n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , 
n17942 , n17944 , n17945 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , 
n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , 
n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , 
n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17982 , n17983 , n17984 , 
n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , 
n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18003 , n18004 , n18005 , n18006 , 
n18007 , n18008 , n18009 , n18010 , n18011 , n18013 , n18014 , n18015 , n18016 , n18017 , 
n18018 , n18019 , n18020 , n18021 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , 
n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18038 , n18039 , 
n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , 
n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , 
n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , 
n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , 
n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18088 , n18089 , n18090 , 
n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , 
n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , 
n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , 
n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , 
n18132 , n18133 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , 
n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , 
n18153 , n18154 , n18155 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , 
n18164 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18175 , 
n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , 
n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , 
n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18205 , n18206 , n18208 , 
n18209 , n18210 , n18211 , n18212 , n18213 , n18215 , n18216 , n18217 , n18218 , n18219 , 
n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , 
n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , 
n18240 , n18241 , n18242 , n18243 , n18244 , n18246 , n18247 , n18248 , n18249 , n18250 , 
n18251 , n18252 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , 
n18262 , n18263 , n18264 , n18265 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , 
n18273 , n18274 , n18275 , n18276 , n18277 , n18279 , n18280 , n18281 , n18282 , n18283 , 
n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18294 , n18295 , 
n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , 
n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , 
n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , 
n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18335 , n18336 , 
n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , 
n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , 
n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , 
n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18377 , 
n18378 , n18379 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18390 , 
n18392 , n18393 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18402 , n18403 , 
n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , 
n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18424 , 
n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , 
n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , 
n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18453 , n18454 , n18455 , n18456 , 
n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , 
n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , 
n18477 , n18478 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , 
n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , 
n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18508 , 
n18509 , n18511 , n18512 , n18513 , n18514 , n18515 , n18517 , n18520 , n18521 , n18522 , 
n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , 
n18533 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , 
n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18552 , n18553 , n18554 , 
n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , 
n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , 
n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18583 , n18584 , n18585 , 
n18586 , n18587 , n18588 , n18589 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , 
n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , 
n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , 
n18617 , n18618 , n18619 , n18620 , n18622 , n18623 , n18624 , n18625 , n18626 , n18628 , 
n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , 
n18641 , n18642 , n18643 , n18644 , n18646 , n18648 , n18649 , n18650 , n18651 , n18652 , 
n18653 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , 
n18664 , n18665 , n18666 , n18668 , n18669 , n18670 , n18671 , n18673 , n18674 , n18675 , 
n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , 
n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , 
n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , 
n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , 
n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , 
n18726 , n18727 , n18728 , n18729 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , 
n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , 
n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , 
n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , 
n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , 
n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , 
n18787 , n18788 , n18789 , n18790 , n18791 , n18793 , n18794 , n18795 , n18796 , n18797 , 
n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , 
n18808 , n18809 , n18811 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , 
n18820 , n18821 , n18822 , n18823 , n18824 , n18826 , n18827 , n18828 , n18829 , n18830 , 
n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , 
n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18851 , 
n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , 
n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , 
n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , 
n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , 
n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , 
n18902 , n18904 , n18905 , n18906 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , 
n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , 
n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , 
n18934 , n18935 , n18936 , n18937 , n18938 , n18940 , n18941 , n18942 , n18943 , n18944 , 
n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , 
n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , 
n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , 
n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , 
n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18994 , n18995 , n18996 , 
n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , 
n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , 
n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19027 , 
n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19036 , n19037 , n19038 , 
n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , 
n19049 , n19050 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , 
n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19067 , n19068 , n19069 , n19070 , 
n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , 
n19081 , n19082 , n19083 , n19084 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , 
n19093 , n19094 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , 
n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19111 , n19112 , n19113 , n19114 , 
n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , 
n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19133 , n19134 , n19135 , 
n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , 
n19147 , n19148 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , 
n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , 
n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , 
n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , 
n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , 
n19198 , n19199 , n19200 , n19201 , n19203 , n19204 , n19206 , n19208 , n19209 , n19210 , 
n19212 , n19213 , n19214 , n19215 , n19216 , n19218 , n19219 , n19220 , n19222 , n19223 , 
n19224 , n19225 , n19226 , n19227 , n19228 , n19230 , n19232 , n19233 , n19234 , n19236 , 
n19237 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , 
n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19256 , n19257 , n19258 , 
n19259 , n19260 , n19262 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , 
n19272 , n19273 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , 
n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , 
n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19301 , n19302 , n19303 , 
n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , 
n19314 , n19315 , n19316 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , 
n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , 
n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , 
n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , 
n19355 , n19357 , n19358 , n19359 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , 
n19367 , n19368 , n19369 , n19370 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , 
n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , 
n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , 
n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19406 , n19407 , n19408 , 
n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , 
n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19426 , n19427 , n19428 , n19429 , 
n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
n19450 , n19451 , n19454 , n19455 , n19456 , n19457 , n19458 , n19460 , n19461 , n19462 , 
n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , 
n19473 , n19474 , n19475 , n19476 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , 
n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , 
n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , 
n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , 
n19514 , n19515 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , 
n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , 
n19535 , n19536 , n19537 , n19539 , n19540 , n19541 , n19543 , n19544 , n19545 , n19547 , 
n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , 
n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , 
n19568 , n19569 , n19570 , n19571 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , 
n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , 
n19590 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , 
n19602 , n19603 , n19605 , n19606 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , 
n19614 , n19616 , n19617 , n19618 , n19619 , n19621 , n19622 , n19623 , n19624 , n19625 , 
n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19633 , n19634 , n19635 , n19636 , 
n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , 
n19647 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , 
n19658 , n19659 , n19660 , n19661 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , 
n19669 , n19670 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , 
n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , 
n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , 
n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , 
n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , 
n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , 
n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , 
n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , 
n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19760 , n19761 , 
n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , 
n19772 , n19773 , n19774 , n19775 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , 
n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , 
n19793 , n19794 , n19795 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , 
n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , 
n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19824 , 
n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , 
n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , 
n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , 
n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , 
n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , 
n19875 , n19876 , n19877 , n19878 , n19879 , n19881 , n19882 , n19883 , n19884 , n19885 , 
n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , 
n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , 
n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , 
n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19924 , n19927 , n19928 , 
n19929 , n19930 , n19931 , n19932 , n19933 , n19935 , n19936 , n19937 , n19938 , n19939 , 
n19940 , n19941 , n19942 , n19944 , n19945 , n19946 , n19947 , n19948 , n19950 , n19951 , 
n19952 , n19953 , n19954 , n19955 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , 
n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , 
n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19981 , n19982 , n19983 , 
n19984 , n19985 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , 
n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , 
n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , 
n20015 , n20016 , n20017 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , 
n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20033 , n20034 , n20035 , n20036 , 
n20037 , n20039 , n20040 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , 
n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , 
n20059 , n20060 , n20061 , n20062 , n20064 , n20066 , n20067 , n20068 , n20069 , n20070 , 
n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20081 , 
n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , 
n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , 
n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , 
n20112 , n20113 , n20114 , n20115 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , 
n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , 
n20133 , n20134 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , 
n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , 
n20154 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , 
n20165 , n20166 , n20167 , n20168 , n20169 , n20171 , n20172 , n20173 , n20174 , n20176 , 
n20177 , n20178 , n20179 , n20180 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , 
n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , 
n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , 
n20209 , n20211 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , 
n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20232 , 
n20233 , n20234 , n20235 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , 
n20244 , n20245 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , 
n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20263 , n20264 , n20265 , 
n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , 
n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , 
n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , 
n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , 
n20306 , n20307 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , 
n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , 
n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , 
n20337 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , 
n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , 
n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20366 , n20367 , n20368 , 
n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , 
n20391 , n20392 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20401 , n20402 , 
n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20411 , n20412 , n20413 , 
n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , 
n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , 
n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20443 , n20444 , 
n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20454 , n20455 , 
n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , 
n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , 
n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20487 , 
n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20496 , n20497 , n20498 , 
n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20508 , n20509 , 
n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , 
n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , 
n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , 
n20541 , n20542 , n20543 , n20544 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , 
n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20561 , n20562 , 
n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , 
n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , 
n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20590 , n20591 , n20592 , n20595 , 
n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , 
n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , 
n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , 
n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20633 , n20634 , n20635 , n20636 , 
n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , 
n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , 
n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20666 , n20667 , n20668 , 
n20669 , n20670 , n20671 , n20672 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , 
n20680 , n20681 , n20682 , n20683 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , 
n20691 , n20692 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , 
n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , 
n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , 
n20722 , n20723 , n20724 , n20725 , n20726 , n20728 , n20729 , n20730 , n20731 , n20732 , 
n20733 , n20734 , n20735 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , 
n20744 , n20745 , n20746 , n20747 , n20748 , n20750 , n20751 , n20752 , n20754 , n20755 , 
n20756 , n20757 , n20758 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , 
n20767 , n20769 , n20770 , n20771 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , 
n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , 
n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , 
n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20809 , n20810 , n20811 , n20813 , 
n20814 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , 
n20826 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , 
n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , 
n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , 
n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , 
n20867 , n20868 , n20869 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , 
n20878 , n20879 , n20880 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , 
n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , 
n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20906 , n20907 , n20908 , n20909 , 
n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , 
n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20930 , 
n20932 , n20933 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , 
n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , 
n20953 , n20954 , n20955 , n20956 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , 
n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , 
n20974 , n20975 , n20977 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , 
n20986 , n20987 , n20988 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , 
n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , 
n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21014 , n21015 , n21016 , n21017 , 
n21018 , n21019 , n21020 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , 
n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , 
n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , 
n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , 
n21059 , n21060 , n21061 , n21062 , n21063 , n21065 , n21066 , n21067 , n21068 , n21069 , 
n21070 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , 
n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , 
n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , 
n21101 , n21102 , n21103 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , 
n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , 
n21123 , n21124 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , 
n21134 , n21135 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , 
n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , 
n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , 
n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , 
n21175 , n21176 , n21178 , n21179 , n21181 , n21182 , n21183 , n21184 , n21187 , n21188 , 
n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , 
n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , 
n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , 
n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , 
n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , 
n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , 
n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , 
n21260 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , 
n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , 
n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , 
n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21300 , n21302 , 
n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , 
n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , 
n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , 
n21334 , n21335 , n21336 , n21337 , n21338 , n21340 , n21341 , n21342 , n21344 , n21345 , 
n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , 
n21357 , n21358 , n21360 , n21361 , n21363 , n21364 , n21366 , n21367 , n21368 , n21369 , 
n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , 
n21380 , n21381 , n21382 , n21383 , n21384 , n21386 , n21387 , n21388 , n21390 , n21391 , 
n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , 
n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , 
n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21422 , n21423 , n21424 , 
n21425 , n21426 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , 
n21436 , n21437 , n21438 , n21439 , n21441 , n21442 , n21443 , n21445 , n21446 , n21447 , 
n21448 , n21449 , n21450 , n21451 , n21452 , n21454 , n21456 , n21457 , n21459 , n21460 , 
n21461 , n21462 , n21463 , n21464 , n21465 , n21467 , n21468 , n21469 , n21471 , n21472 , 
n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , 
n21483 , n21484 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21494 , 
n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , 
n21505 , n21506 , n21507 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , 
n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , 
n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , 
n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21546 , 
n21547 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , 
n21559 , n21560 , n21561 , n21562 , n21564 , n21565 , n21566 , n21567 , n21568 , n21570 , 
n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , 
n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , 
n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21598 , n21599 , n21600 , n21601 , 
n21602 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , 
n21613 , n21614 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , 
n21624 , n21625 , n21626 , n21627 , n21629 , n21630 , n21631 , n21633 , n21634 , n21635 , 
n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , 
n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21654 , n21656 , n21657 , 
n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , 
n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , 
n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21687 , n21689 , 
n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , 
n21700 , n21701 , n21703 , n21704 , n21705 , n21707 , n21709 , n21710 , n21711 , n21712 , 
n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21723 , 
n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , 
n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , 
n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , 
n21754 , n21755 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , 
n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21772 , n21773 , n21774 , n21775 , 
n21776 , n21777 , n21778 , n21779 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , 
n21788 , n21789 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , 
n21799 , n21800 , n21802 , n21803 , n21804 , n21805 , n21807 , n21809 , n21810 , n21811 , 
n21812 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , 
n21823 , n21824 , n21825 , n21826 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , 
n21834 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , 
n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , 
n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21863 , n21865 , n21866 , 
n21867 , n21868 , n21869 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , 
n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , 
n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , 
n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , 
n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21919 , 
n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , 
n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , 
n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , 
n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , 
n21961 , n21962 , n21964 , n21965 , n21967 , n21968 , n21969 , n21971 , n21972 , n21973 , 
n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , 
n21984 , n21985 , n21986 , n21987 , n21988 , n21990 , n21991 , n21992 , n21993 , n21994 , 
n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , 
n22005 , n22006 , n22007 , n22008 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , 
n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , 
n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , 
n22036 , n22037 , n22038 , n22039 , n22041 , n22042 , n22043 , n22044 , n22046 , n22047 , 
n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , 
n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , 
n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22076 , n22077 , n22078 , 
n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , 
n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , 
n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , 
n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22117 , n22119 , n22120 , 
n22122 , n22123 , n22124 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , 
n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , 
n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , 
n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , 
n22163 , n22165 , n22166 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , 
n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22186 , 
n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , 
n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22206 , n22208 , 
n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22219 , 
n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , 
n22230 , n22231 , n22232 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , 
n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , 
n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22258 , n22259 , n22260 , n22261 , 
n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22271 , n22272 , 
n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , 
n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , 
n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , 
n22303 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , 
n22315 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , 
n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , 
n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , 
n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , 
n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , 
n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , 
n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , 
n22387 , n22389 , n22390 , n22391 , n22392 , n22394 , n22395 , n22396 , n22397 , n22398 , 
n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , 
n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , 
n22419 , n22420 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , 
n22432 , n22433 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , 
n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22452 , n22453 , n22454 , 
n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , 
n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , 
n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , 
n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , 
n22495 , n22496 , n22497 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , 
n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22513 , n22514 , n22515 , n22516 , 
n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , 
n22527 , n22528 , n22529 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , 
n22538 , n22539 , n22540 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , 
n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , 
n22561 , n22562 , n22563 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , 
n22572 , n22573 , n22574 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , 
n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , 
n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22601 , n22602 , n22604 , 
n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , 
n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , 
n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22634 , n22635 , 
n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , 
n22646 , n22647 , n22648 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , 
n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22668 , n22669 , 
n22670 , n22671 , n22672 , n22673 , n22674 , n22676 , n22677 , n22679 , n22680 , n22681 , 
n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , 
n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22703 , 
n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22714 , 
n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , 
n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , 
n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , 
n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , 
n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , 
n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22774 , n22775 , n22776 , 
n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , 
n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , 
n22797 , n22798 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , 
n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , 
n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , 
n22828 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , 
n22840 , n22841 , n22842 , n22843 , n22844 , n22846 , n22847 , n22848 , n22849 , n22850 , 
n22851 , n22852 , n22853 , n22854 , n22855 , n22857 , n22858 , n22859 , n22860 , n22861 , 
n22862 , n22863 , n22865 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , 
n22875 , n22876 , n22877 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , 
n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , 
n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , 
n22907 , n22908 , n22910 , n22911 , n22912 , n22914 , n22915 , n22916 , n22918 , n22919 , 
n22921 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22930 , n22931 , n22932 , 
n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , 
n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , 
n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22961 , n22963 , n22964 , 
n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , 
n22975 , n22976 , n22977 , n22978 , n22980 , n22981 , n22982 , n22983 , n22984 , n22986 , 
n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , 
n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , 
n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , 
n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23024 , n23025 , n23026 , n23027 , 
n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , 
n23038 , n23039 , n23041 , n23042 , n23044 , n23045 , n23048 , n23049 , n23050 , n23051 , 
n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , 
n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23072 , n23073 , 
n23074 , n23075 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , 
n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , 
n23095 , n23096 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , 
n23106 , n23107 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23116 , n23117 , 
n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , 
n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , 
n23138 , n23139 , n23140 , n23141 , n23142 , n23146 , n23147 , n23148 , n23149 , n23150 , 
n23151 , n23152 , n23153 , n23154 , n23155 , n23157 , n23158 , n23159 , n23160 , n23161 , 
n23162 , n23163 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , 
n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , 
n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , 
n23194 , n23196 , n23197 , n23198 , n23200 , n23201 , n23202 , n23203 , n23205 , n23206 , 
n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , 
n23217 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , 
n23228 , n23229 , n23230 , n23231 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , 
n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , 
n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , 
n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , 
n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , 
n23279 , n23280 , n23281 , n23283 , n23284 , n23285 , n23286 , n23287 , n23289 , n23290 , 
n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , 
n23301 , n23302 , n23303 , n23305 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , 
n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23321 , n23322 , n23323 , 
n23324 , n23325 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , 
n23335 , n23337 , n23338 , n23339 , n23340 , n23341 , n23343 , n23344 , n23345 , n23346 , 
n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , 
n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , 
n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23376 , n23377 , n23378 , 
n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , 
n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , 
n23399 , n23401 , n23402 , n23404 , n23405 , n23408 , n23409 , n23410 , n23411 , n23412 , 
n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23420 , n23421 , n23422 , n23423 , 
n23424 , n23425 , n23426 , n23427 , n23428 , n23430 , n23432 , n23433 , n23434 , n23435 , 
n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , 
n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , 
n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23465 , n23466 , 
n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , 
n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , 
n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , 
n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , 
n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , 
n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , 
n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , 
n23537 , n23538 , n23539 , n23541 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , 
n23549 , n23550 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23559 , n23562 , 
n23563 , n23564 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , 
n23574 , n23575 , n23576 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , 
n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , 
n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , 
n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , 
n23615 , n23616 , n23617 , n23618 , n23619 , n23621 , n23622 , n23623 , n23624 , n23625 , 
n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , 
n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23644 , n23645 , n23646 , 
n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23656 , n23657 , 
n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , 
n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , 
n23678 , n23679 , n23680 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , 
n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , 
n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , 
n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , 
n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , 
n23729 , n23730 , n23731 , n23732 , n23733 , n23735 , n23736 , n23737 , n23738 , n23739 , 
n23740 , n23741 , n23742 , n23743 , n23745 , n23746 , n23747 , n23748 , n23750 , n23751 , 
n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , 
n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23772 , n23773 , 
n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , 
n23784 , n23785 , n23786 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , 
n23795 , n23796 , n23797 , n23798 , n23799 , n23801 , n23802 , n23803 , n23804 , n23805 , 
n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , 
n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23825 , n23826 , 
n23827 , n23828 , n23829 , n23830 , n23831 , n23833 , n23834 , n23836 , n23837 , n23839 , 
n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , 
n23850 , n23851 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
n23901 , n23902 , n23903 , n23904 , n23905 , n23907 , n23908 , n23909 , n23910 , n23911 , 
n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , 
n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , 
n23933 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , 
n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , 
n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23961 , n23962 , n23963 , n23964 , 
n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , 
n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , 
n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , 
n23995 , n23996 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , 
n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , 
n24016 , n24017 , n24018 , n24019 , n24020 , n24023 , n24024 , n24025 , n24026 , n24027 , 
n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , 
n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24048 , 
n24049 , n24050 , n24051 , n24052 , n24054 , n24055 , n24057 , n24058 , n24059 , n24060 , 
n24061 , n24062 , n24063 , n24064 , n24065 , n24067 , n24068 , n24069 , n24070 , n24071 , 
n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , 
n24082 , n24083 , n24084 , n24085 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , 
n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24101 , n24102 , n24103 , 
n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , 
n24115 , n24116 , n24117 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , 
n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24133 , n24134 , n24135 , n24136 , 
n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24145 , n24146 , n24147 , n24148 , 
n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , 
n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , 
n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , 
n24180 , n24181 , n24182 , n24183 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
n24211 , n24212 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , 
n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , 
n24233 , n24234 , n24235 , n24236 , n24237 , n24239 , n24240 , n24241 , n24242 , n24243 , 
n24244 , n24245 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , 
n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , 
n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , 
n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24284 , n24285 , 
n24286 , n24287 , n24288 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , 
n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24305 , n24306 , n24307 , 
n24308 , n24309 , n24310 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , 
n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , 
n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24339 , 
n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , 
n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24378 , n24379 , n24380 , n24381 , 
n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , 
n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24399 , n24400 , n24401 , n24402 , 
n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , 
n24413 , n24414 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , 
n24424 , n24425 , n24426 , n24427 , n24428 , n24430 , n24431 , n24432 , n24433 , n24434 , 
n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , 
n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , 
n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24465 , n24466 , 
n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24474 , n24475 , n24476 , n24477 , 
n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , 
n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , 
n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , 
n24509 , n24510 , n24511 , n24513 , n24514 , n24516 , n24517 , n24518 , n24519 , n24520 , 
n24521 , n24523 , n24524 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , 
n24534 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , 
n24545 , n24546 , n24547 , n24548 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , 
n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , 
n24566 , n24567 , n24568 , n24570 , n24571 , n24572 , n24573 , n24574 , n24576 , n24577 , 
n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24587 , n24588 , n24589 , 
n24590 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24629 , n24630 , n24631 , 
n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , 
n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24649 , n24650 , n24651 , n24652 , 
n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , 
n24663 , n24664 , n24665 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , 
n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , 
n24684 , n24685 , n24686 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , 
n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , 
n24705 , n24706 , n24707 , n24709 , n24710 , n24711 , n24713 , n24714 , n24715 , n24716 , 
n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24745 , n24746 , n24747 , 
n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , 
n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24768 , 
n24769 , n24771 , n24772 , n24773 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24790 , n24791 , 
n24792 , n24793 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , 
n24805 , n24806 , n24809 , n24810 , n24812 , n24813 , n24814 , n24815 , n24816 , n24818 , 
n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , 
n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24838 , n24839 , 
n24840 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
n24881 , n24882 , n24883 , n24884 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , 
n24893 , n24894 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , 
n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , 
n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , 
n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , 
n24934 , n24935 , n24936 , n24938 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , 
n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , 
n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , 
n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , 
n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , 
n24987 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , 
n24998 , n25000 , n25001 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , 
n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , 
n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , 
n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , 
n25040 , n25041 , n25042 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , 
n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25090 , n25091 , 
n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , 
n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , 
n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , 
n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , 
n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , 
n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , 
n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , 
n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25173 , n25174 , n25175 , 
n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , 
n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25194 , n25195 , n25196 , 
n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , 
n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , 
n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , 
n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25236 , n25237 , 
n25238 , n25239 , n25240 , n25241 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
n25249 , n25250 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , 
n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , 
n25270 , n25271 , n25272 , n25274 , n25275 , n25277 , n25278 , n25279 , n25280 , n25281 , 
n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25292 , 
n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , 
n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25311 , n25312 , n25313 , 
n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , 
n25324 , n25325 , n25326 , n25327 , n25328 , n25330 , n25331 , n25332 , n25333 , n25335 , 
n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , 
n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , 
n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , 
n25366 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , 
n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , 
n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25397 , 
n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , 
n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , 
n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , 
n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , 
n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , 
n25449 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , 
n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , 
n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , 
n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25488 , n25489 , n25490 , 
n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , 
n25501 , n25503 , n25504 , n25505 , n25506 , n25507 , n25510 , n25511 , n25512 , n25513 , 
n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , 
n25524 , n25525 , n25526 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , 
n25535 , n25536 , n25537 , n25538 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , 
n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , 
n25556 , n25557 , n25558 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , 
n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , 
n25577 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25587 , n25588 , n25589 , 
n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , 
n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , 
n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , 
n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , 
n25630 , n25631 , n25632 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , 
n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , 
n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , 
n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , 
n25672 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , 
n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , 
n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25700 , n25701 , n25702 , n25703 , 
n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , 
n25714 , n25715 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25743 , n25744 , n25745 , n25746 , 
n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , 
n25757 , n25759 , n25761 , n25762 , n25763 , n25765 , n25766 , n25767 , n25768 , n25769 , 
n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , 
n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , 
n25791 , n25792 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , 
n25802 , n25803 , n25804 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , 
n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , 
n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , 
n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , 
n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , 
n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , 
n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25871 , n25872 , n25873 , n25874 , 
n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
n25885 , n25886 , n25887 , n25888 , n25890 , n25892 , n25893 , n25894 , n25895 , n25896 , 
n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , 
n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , 
n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , 
n25927 , n25928 , n25929 , n25931 , n25932 , n25933 , n25935 , n25936 , n25937 , n25938 , 
n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25946 , n25947 , n25948 , n25949 , 
n25950 , n25951 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , 
n25961 , n25962 , n25964 , n25965 , n25966 , n25967 , n25969 , n25970 , n25971 , n25972 , 
n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , 
n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25990 , n25992 , n25993 , n25994 , 
n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26003 , n26005 , n26006 , n26008 , 
n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , 
n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , 
n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , 
n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , 
n26049 , n26050 , n26051 , n26053 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , 
n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , 
n26071 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , 
n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26091 , n26092 , n26093 , 
n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26104 , n26105 , 
n26106 , n26107 , n26109 , n26110 , n26111 , n26112 , n26113 , n26116 , n26117 , n26118 , 
n26119 , n26120 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , 
n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , 
n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26150 , 
n26151 , n26152 , n26154 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , 
n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , 
n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , 
n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26192 , n26193 , n26194 , 
n26195 , n26196 , n26198 , n26199 , n26200 , n26201 , n26202 , n26204 , n26205 , n26206 , 
n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , 
n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , 
n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , 
n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , 
n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , 
n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , 
n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , 
n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , 
n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , 
n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26307 , 
n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , 
n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , 
n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26336 , n26337 , n26338 , 
n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , 
n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , 
n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26416 , n26417 , n26418 , n26419 , 
n26420 , n26421 , n26422 , n26423 , n26424 , n26426 , n26427 , n26428 , n26429 , n26430 , 
n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , 
n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26448 , n26449 , n26450 , n26451 , 
n26452 , n26453 , n26454 , n26455 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , 
n26463 , n26464 , n26465 , n26467 , n26468 , n26469 , n26471 , n26472 , n26473 , n26474 , 
n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
n26505 , n26506 , n26507 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , 
n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , 
n26527 , n26528 , n26529 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , 
n26538 , n26539 , n26540 , n26542 , n26543 , n26544 , n26545 , n26546 , n26548 , n26549 , 
n26550 , n26551 , n26552 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , 
n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , 
n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26580 , n26581 , n26582 , 
n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , 
n26593 , n26594 , n26595 , n26596 , n26597 , n26599 , n26600 , n26601 , n26602 , n26603 , 
n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , 
n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , 
n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , 
n26634 , n26635 , n26637 , n26638 , n26639 , n26640 , n26641 , n26643 , n26644 , n26645 , 
n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , 
n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26666 , 
n26667 , n26668 , n26669 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , 
n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , 
n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26695 , n26696 , n26697 , n26698 , 
n26699 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , 
n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , 
n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26730 , 
n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , 
n26742 , n26743 , n26744 , n26745 , n26746 , n26748 , n26749 , n26750 , n26751 , n26752 , 
n26753 , n26754 , n26755 , n26756 , n26757 , n26759 , n26760 , n26761 , n26762 , n26763 , 
n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
n26775 , n26776 , n26777 , n26779 , n26780 , n26782 , n26783 , n26784 , n26787 , n26788 , 
n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , 
n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , 
n26809 , n26810 , n26811 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , 
n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , 
n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26838 , n26840 , n26841 , 
n26842 , n26843 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , 
n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , 
n26864 , n26865 , n26866 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
n26875 , n26876 , n26877 , n26878 , n26879 , n26881 , n26882 , n26883 , n26884 , n26886 , 
n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26895 , n26896 , n26897 , 
n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , 
n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , 
n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , 
n26930 , n26931 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26941 , 
n26942 , n26943 , n26944 , n26945 , n26946 , n26948 , n26949 , n26950 , n26951 , n26952 , 
n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26962 , n26963 , n26965 , 
n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26975 , n26976 , 
n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , 
n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26997 , 
n26998 , n26999 , n27000 , n27001 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , 
n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , 
n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
n27029 , n27030 , n27031 , n27032 , n27033 , n27035 , n27036 , n27037 , n27038 , n27039 , 
n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , 
n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27057 , n27058 , n27059 , n27060 , 
n27061 , n27062 , n27063 , n27065 , n27066 , n27067 , n27068 , n27069 , n27071 , n27072 , 
n27073 , n27074 , n27075 , n27076 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , 
n27084 , n27086 , n27087 , n27088 , n27089 , n27091 , n27092 , n27093 , n27094 , n27096 , 
n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , 
n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , 
n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27127 , 
n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27135 , n27136 , n27137 , n27138 , 
n27139 , n27140 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , 
n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , 
n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , 
n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , 
n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , 
n27191 , n27192 , n27193 , n27194 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , 
n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27212 , 
n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , 
n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27234 , 
n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27253 , n27255 , n27256 , 
n27257 , n27258 , n27259 , n27260 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , 
n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , 
n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , 
n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , 
n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27306 , n27307 , n27308 , 
n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27316 , n27317 , n27319 , n27320 , 
n27321 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , 
n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , 
n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , 
n27352 , n27353 , n27357 , n27358 , n27359 , n27360 , n27362 , n27363 , n27364 , n27365 , 
n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , 
n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , 
n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , 
n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , 
n27407 , n27408 , n27409 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , 
n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , 
n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , 
n27438 , n27439 , n27440 , n27441 , n27442 , n27444 , n27445 , n27446 , n27447 , n27448 , 
n27449 , n27450 , n27451 , n27452 , n27454 , n27455 , n27457 , n27458 , n27459 , n27460 , 
n27461 , n27462 , n27463 , n27465 , n27466 , n27468 , n27469 , n27470 , n27471 , n27473 , 
n27474 , n27475 , n27476 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , 
n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27493 , n27494 , n27495 , 
n27496 , n27497 , n27498 , n27499 , n27500 , n27503 , n27504 , n27505 , n27507 , n27509 , 
n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , 
n27520 , n27521 , n27522 , n27523 , n27525 , n27526 , n27527 , n27529 , n27530 , n27531 , 
n27532 , n27533 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , 
n27543 , n27544 , n27545 , n27546 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , 
n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , 
n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27573 , n27574 , n27575 , n27576 , 
n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , 
n27587 , n27588 , n27589 , n27590 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , 
n27598 , n27599 , n27600 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , 
n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , 
n27619 , n27620 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , 
n27630 , n27631 , n27633 , n27634 , n27635 , n27637 , n27638 , n27640 , n27641 , n27642 , 
n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , 
n27653 , n27654 , n27655 , n27656 , n27657 , n27659 , n27660 , n27661 , n27662 , n27663 , 
n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , 
n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , 
n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , 
n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , 
n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27714 , 
n27715 , n27716 , n27717 , n27718 , n27719 , n27721 , n27722 , n27723 , n27724 , n27725 , 
n27726 , n27727 , n27728 , n27729 , n27731 , n27732 , n27733 , n27734 , n27735 , n27737 , 
n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , 
n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , 
n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , 
n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , 
n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , 
n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , 
n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27806 , n27807 , n27808 , 
n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , 
n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , 
n27830 , n27831 , n27832 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , 
n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27849 , n27850 , n27851 , 
n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , 
n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , 
n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , 
n27884 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , 
n27897 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , 
n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , 
n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , 
n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , 
n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , 
n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , 
n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , 
n27969 , n27970 , n27971 , n27972 , n27973 , n27975 , n27976 , n27977 , n27978 , n27979 , 
n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , 
n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , 
n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28007 , n28008 , n28009 , n28010 , 
n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , 
n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , 
n28031 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , 
n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , 
n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , 
n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , 
n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28082 , 
n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , 
n28093 , n28094 , n28095 , n28096 , n28097 , n28099 , n28100 , n28101 , n28102 , n28103 , 
n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28114 , 
n28115 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28125 , n28126 , 
n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , 
n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28147 , n28148 , 
n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28159 , 
n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , 
n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , 
n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28189 , n28190 , n28191 , 
n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , 
n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , 
n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , 
n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , 
n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , 
n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , 
n28252 , n28253 , n28254 , n28255 , n28256 , n28258 , n28259 , n28260 , n28261 , n28262 , 
n28263 , n28264 , n28265 , n28266 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , 
n28274 , n28275 , n28276 , n28277 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , 
n28285 , n28286 , n28287 , n28288 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , 
n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28306 , 
n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , 
n28317 , n28318 , n28319 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , 
n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28338 , 
n28339 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , 
n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , 
n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , 
n28370 , n28371 , n28372 , n28373 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , 
n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , 
n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28398 , n28400 , n28401 , n28403 , 
n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , 
n28414 , n28415 , n28418 , n28419 , n28420 , n28421 , n28423 , n28424 , n28425 , n28426 , 
n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28434 , n28435 , n28436 , n28437 , 
n28438 , n28439 , n28440 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , 
n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , 
n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , 
n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , 
n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , 
n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , 
n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , 
n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28518 , n28519 , 
n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , 
n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28538 , n28539 , n28540 , 
n28541 , n28542 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , 
n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28563 , 
n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , 
n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , 
n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , 
n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28605 , 
n28607 , n28608 , n28610 , n28611 , n28612 , n28614 , n28615 , n28616 , n28617 , n28618 , 
n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , 
n28629 , n28630 , n28631 , n28632 , n28633 , n28635 , n28637 , n28639 , n28640 , n28641 , 
n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , 
n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , 
n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28671 , n28672 , 
n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28682 , n28683 , 
n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , 
n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28704 , 
n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , 
n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , 
n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28735 , 
n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , 
n28746 , n28747 , n28748 , n28749 , n28751 , n28752 , n28753 , n28755 , n28756 , n28757 , 
n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , 
n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , 
n28778 , n28779 , n28780 , n28782 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , 
n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , 
n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , 
n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , 
n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28829 , n28830 , 
n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , 
n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , 
n28851 , n28853 , n28854 , n28855 , n28857 , n28858 , n28859 , n28861 , n28862 , n28863 , 
n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , 
n28874 , n28875 , n28876 , n28877 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , 
n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , 
n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , 
n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , 
n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , 
n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28944 , n28945 , 
n28946 , n28947 , n28948 , n28949 , n28950 , n28953 , n28954 , n28955 , n28956 , n28958 , 
n28959 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , 
n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , 
n28980 , n28981 , n28982 , n28984 , n28985 , n28986 , n28987 , n28988 , n28990 , n28991 , 
n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29002 , 
n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , 
n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , 
n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29032 , n29033 , n29034 , 
n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , 
n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , 
n29055 , n29056 , n29057 , n29058 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , 
n29066 , n29067 , n29068 , n29069 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , 
n29077 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , 
n29088 , n29089 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , 
n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , 
n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , 
n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , 
n29129 , n29130 , n29131 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , 
n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , 
n29150 , n29151 , n29152 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , 
n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , 
n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , 
n29181 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29190 , n29191 , n29192 , 
n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , 
n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , 
n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , 
n29223 , n29224 , n29225 , n29226 , n29228 , n29230 , n29231 , n29232 , n29233 , n29234 , 
n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , 
n29245 , n29246 , n29247 , n29248 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , 
n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29266 , 
n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , 
n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , 
n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29294 , n29295 , n29296 , n29297 , 
n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29307 , n29308 , 
n29309 , n29310 , n29311 , n29312 , n29313 , n29315 , n29317 , n29318 , n29319 , n29320 , 
n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , 
n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , 
n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , 
n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29361 , 
n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29370 , n29371 , n29372 , 
n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29381 , n29383 , n29384 , 
n29385 , n29386 , n29387 , n29388 , n29389 , n29391 , n29392 , n29393 , n29394 , n29395 , 
n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , 
n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , 
n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , 
n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29438 , 
n29439 , n29440 , n29441 , n29442 , n29443 , n29445 , n29446 , n29448 , n29449 , n29451 , 
n29452 , n29453 , n29454 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , 
n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29472 , n29473 , n29474 , 
n29475 , n29476 , n29477 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , 
n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , 
n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , 
n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , 
n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , 
n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , 
n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , 
n29546 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , 
n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29567 , 
n29568 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , 
n29579 , n29580 , n29581 , n29582 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , 
n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , 
n29600 , n29601 , n29602 , n29603 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , 
n29611 , n29612 , n29613 , n29614 , n29616 , n29617 , n29618 , n29620 , n29621 , n29622 , 
n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , 
n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , 
n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29651 , n29652 , n29653 , n29654 , 
n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29663 , n29664 , n29665 , 
n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29678 , n29679 , 
n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , 
n29690 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , 
n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29712 , n29713 , 
n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29721 , n29722 , n29723 , n29724 , 
n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , 
n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , 
n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , 
n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29765 , n29766 , 
n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , 
n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , 
n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , 
n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29805 , n29806 , n29807 , 
n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , 
n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , 
n29829 , n29830 , n29831 , n29832 , n29834 , n29835 , n29836 , n29837 , n29839 , n29840 , 
n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , 
n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , 
n29861 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , 
n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29879 , n29880 , n29881 , n29882 , 
n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , 
n29894 , n29895 , n29896 , n29898 , n29899 , n29900 , n29901 , n29903 , n29904 , n29905 , 
n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , 
n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , 
n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29934 , n29935 , n29936 , 
n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , 
n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , 
n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , 
n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29975 , n29976 , n29977 , 
n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , 
n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29997 , n29998 , n29999 , 
n30000 , n30001 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30010 , n30011 , 
n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , 
n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , 
n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , 
n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , 
n30053 , n30054 , n30055 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , 
n30064 , n30065 , n30066 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , 
n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , 
n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , 
n30095 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , 
n30106 , n30107 , n30108 , n30109 , n30110 , n30112 , n30113 , n30114 , n30115 , n30116 , 
n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , 
n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , 
n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , 
n30147 , n30148 , n30149 , n30151 , n30152 , n30154 , n30155 , n30156 , n30157 , n30159 , 
n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30168 , n30169 , n30171 , 
n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , 
n30183 , n30184 , n30185 , n30186 , n30187 , n30189 , n30190 , n30191 , n30192 , n30193 , 
n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30202 , n30203 , n30204 , 
n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , 
n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , 
n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , 
n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , 
n30246 , n30247 , n30248 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , 
n30258 , n30259 , n30261 , n30262 , n30263 , n30264 , n30265 , n30267 , n30268 , n30270 , 
n30271 , n30272 , n30273 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , 
n30283 , n30284 , n30285 , n30286 , n30288 , n30290 , n30291 , n30292 , n30293 , n30294 , 
n30295 , n30296 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , 
n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , 
n30316 , n30317 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30327 , 
n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , 
n30338 , n30339 , n30340 , n30341 , n30342 , n30344 , n30345 , n30346 , n30347 , n30348 , 
n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , 
n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , 
n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , 
n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , 
n30389 , n30390 , n30391 , n30392 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , 
n30400 , n30401 , n30402 , n30403 , n30404 , n30406 , n30407 , n30408 , n30409 , n30410 , 
n30412 , n30413 , n30414 , n30415 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , 
n30423 , n30424 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30433 , n30434 , 
n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , 
n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , 
n30456 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , 
n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , 
n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , 
n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , 
n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30506 , n30507 , n30508 , 
n30509 , n30510 , n30511 , n30512 , n30513 , n30515 , n30516 , n30517 , n30518 , n30519 , 
n30520 , n30521 , n30522 , n30523 , n30524 , n30526 , n30527 , n30528 , n30530 , n30531 , 
n30532 , n30533 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , 
n30544 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , 
n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30563 , n30564 , n30565 , 
n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , 
n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , 
n30588 , n30589 , n30590 , n30591 , n30592 , n30594 , n30595 , n30596 , n30597 , n30598 , 
n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , 
n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , 
n30619 , n30620 , n30621 , n30622 , n30623 , n30626 , n30627 , n30628 , n30629 , n30630 , 
n30631 , n30632 , n30633 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , 
n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , 
n30652 , n30653 , n30654 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , 
n30663 , n30665 , n30666 , n30667 , n30668 , n30670 , n30671 , n30672 , n30673 , n30674 , 
n30675 , n30676 , n30677 , n30678 , n30680 , n30681 , n30682 , n30683 , n30684 , n30686 , 
n30687 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , 
n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30707 , n30708 , 
n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , 
n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30728 , n30730 , 
n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , 
n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , 
n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , 
n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30770 , n30771 , 
n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , 
n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30789 , n30790 , n30791 , n30792 , 
n30793 , n30794 , n30795 , n30796 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , 
n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , 
n30816 , n30817 , n30818 , n30819 , n30820 , n30822 , n30823 , n30824 , n30825 , n30826 , 
n30827 , n30828 , n30829 , n30830 , n30832 , n30833 , n30834 , n30835 , n30836 , n30838 , 
n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30847 , n30848 , n30849 , n30850 , 
n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , 
n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , 
n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , 
n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30888 , n30889 , n30890 , n30891 , 
n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , 
n30903 , n30904 , n30905 , n30906 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , 
n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , 
n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , 
n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , 
n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30955 , n30956 , n30957 , n30958 , 
n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , 
n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , 
n30979 , n30980 , n30981 , n30982 , n30983 , n30985 , n30986 , n30987 , n30988 , n30989 , 
n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , 
n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , 
n31010 , n31011 , n31013 , n31014 , n31016 , n31018 , n31020 , n31021 , n31022 , n31023 , 
n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , 
n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , 
n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , 
n31054 , n31056 , n31057 , n31059 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , 
n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31074 , n31075 , n31076 , n31078 , 
n31079 , n31080 , n31081 , n31082 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , 
n31090 , n31091 , n31092 , n31093 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , 
n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31109 , n31110 , n31112 , 
n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , 
n31123 , n31124 , n31125 , n31126 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , 
n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31145 , 
n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , 
n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , 
n31166 , n31167 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , 
n31177 , n31178 , n31179 , n31180 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , 
n31188 , n31190 , n31191 , n31192 , n31193 , n31195 , n31196 , n31198 , n31199 , n31200 , 
n31201 , n31202 , n31203 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , 
n31212 , n31213 , n31214 , n31215 , n31216 , n31218 , n31219 , n31220 , n31222 , n31223 , 
n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , 
n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , 
n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , 
n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31265 , 
n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , 
n31276 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31287 , 
n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , 
n31298 , n31299 , n31300 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , 
n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , 
n31319 , n31320 , n31322 , n31323 , n31324 , n31325 , n31327 , n31328 , n31329 , n31330 , 
n31331 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , 
n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31350 , n31352 , n31353 , 
n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , 
n31364 , n31365 , n31367 , n31368 , n31369 , n31371 , n31372 , n31374 , n31375 , n31376 , 
n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , 
n31387 , n31388 , n31389 , n31391 , n31392 , n31393 , n31394 , n31395 , n31398 , n31399 , 
n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , 
n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , 
n31420 , n31422 , n31423 , n31424 , n31425 , n31427 , n31428 , n31429 , n31430 , n31431 , 
n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , 
n31442 , n31443 , n31444 , n31445 , n31446 , n31449 , n31450 , n31451 , n31452 , n31453 , 
n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , 
n31464 , n31465 , n31467 , n31468 , n31469 , n31471 , n31472 , n31473 , n31474 , n31475 , 
n31476 , n31477 , n31478 , n31479 , n31480 , n31482 , n31483 , n31485 , n31486 , n31487 , 
n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , 
n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31506 , n31507 , n31508 , 
n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , 
n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , 
n31529 , n31530 , n31531 , n31532 , n31533 , n31535 , n31537 , n31538 , n31539 , n31540 , 
n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , 
n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , 
n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31571 , 
n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , 
n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31592 , 
n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , 
n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , 
n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , 
n31623 , n31624 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , 
n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , 
n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31651 , n31652 , n31653 , n31654 , 
n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , 
n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , 
n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , 
n31685 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31694 , n31695 , n31696 , 
n31697 , n31698 , n31699 , n31700 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , 
n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , 
n31718 , n31719 , n31720 , n31721 , n31723 , n31724 , n31726 , n31728 , n31729 , n31730 , 
n31731 , n31732 , n31734 , n31735 , n31737 , n31738 , n31739 , n31740 , n31742 , n31743 , 
n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , 
n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31764 , n31765 , n31766 , 
n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31774 , n31775 , n31776 , n31777 , 
n31778 , n31779 , n31780 , n31781 , n31782 , n31785 , n31786 , n31787 , n31788 , n31790 , 
n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , 
n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , 
n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , 
n31821 , n31822 , n31823 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , 
n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , 
n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31849 , n31850 , n31851 , n31852 , 
n31853 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , 
n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , 
n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , 
n31884 , n31885 , n31886 , n31887 , n31888 , n31890 , n31891 , n31892 , n31893 , n31894 , 
n31895 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , 
n31906 , n31908 , n31909 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , 
n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , 
n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , 
n31938 , n31939 , n31941 , n31942 , n31943 , n31944 , n31946 , n31947 , n31948 , n31949 , 
n31950 , n31951 , n31952 , n31953 , n31954 , n31956 , n31957 , n31958 , n31959 , n31960 , 
n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31971 , 
n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31982 , 
n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31991 , n31992 , n31993 , 
n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , 
n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , 
n32014 , n32015 , n32016 , n32017 , n32019 , n32020 , n32021 , n32022 , n32024 , n32025 , 
n32026 , n32027 , n32028 , n32030 , n32031 , n32032 , n32033 , n32034 ;
    not g0 ( n15827 , n6024 );
    and g1 ( n9764 , n30631 , n24174 );
    not g2 ( n18060 , n4981 );
    and g3 ( n20286 , n2939 , n23040 );
    not g4 ( n29665 , n17531 );
    or g5 ( n8383 , n13195 , n4892 );
    or g6 ( n5467 , n516 , n11608 );
    or g7 ( n861 , n16957 , n23102 );
    xnor g8 ( n689 , n8555 , n22867 );
    xnor g9 ( n23571 , n1746 , n9395 );
    or g10 ( n10256 , n2171 , n7607 );
    not g11 ( n26502 , n19440 );
    xnor g12 ( n20684 , n31880 , n4680 );
    and g13 ( n2609 , n19969 , n31268 );
    not g14 ( n19215 , n24775 );
    and g15 ( n12034 , n22155 , n19391 );
    nor g16 ( n17135 , n30646 , n9194 );
    nor g17 ( n13801 , n7690 , n1397 );
    and g18 ( n11619 , n18874 , n3253 );
    xnor g19 ( n1480 , n19368 , n4286 );
    not g20 ( n27581 , n18768 );
    xnor g21 ( n9244 , n30294 , n6005 );
    not g22 ( n8021 , n19458 );
    not g23 ( n2103 , n14812 );
    nor g24 ( n6851 , n6433 , n29533 );
    xnor g25 ( n8008 , n14701 , n18126 );
    or g26 ( n27418 , n11718 , n1551 );
    not g27 ( n31608 , n25336 );
    xnor g28 ( n26479 , n23744 , n15100 );
    xnor g29 ( n23041 , n20825 , n13494 );
    or g30 ( n5429 , n14046 , n30283 );
    nor g31 ( n10157 , n19425 , n22936 );
    not g32 ( n8457 , n12540 );
    and g33 ( n25852 , n10384 , n4543 );
    and g34 ( n2051 , n12307 , n13617 );
    or g35 ( n25051 , n8660 , n31297 );
    not g36 ( n23163 , n12511 );
    and g37 ( n8766 , n31978 , n1224 );
    or g38 ( n13117 , n6094 , n4874 );
    xnor g39 ( n15742 , n3072 , n14978 );
    or g40 ( n13911 , n13846 , n31898 );
    not g41 ( n7029 , n1084 );
    not g42 ( n26193 , n20164 );
    or g43 ( n17237 , n15644 , n25638 );
    xnor g44 ( n27195 , n8103 , n8953 );
    xor g45 ( n15945 , n4434 , n19350 );
    or g46 ( n5343 , n15552 , n8756 );
    or g47 ( n27399 , n15690 , n25985 );
    or g48 ( n15067 , n20116 , n18604 );
    and g49 ( n32006 , n4079 , n3387 );
    not g50 ( n31798 , n25495 );
    and g51 ( n31644 , n24030 , n25244 );
    or g52 ( n14215 , n13349 , n28698 );
    xnor g53 ( n4760 , n21918 , n6651 );
    nor g54 ( n8608 , n14370 , n17979 );
    not g55 ( n18402 , n15224 );
    xnor g56 ( n21268 , n24377 , n28113 );
    or g57 ( n598 , n30471 , n24388 );
    not g58 ( n4614 , n19534 );
    xnor g59 ( n7426 , n2264 , n12605 );
    nor g60 ( n3847 , n4583 , n30906 );
    nor g61 ( n25483 , n3853 , n27633 );
    and g62 ( n8861 , n9827 , n27741 );
    nor g63 ( n29451 , n9801 , n26725 );
    or g64 ( n31014 , n6874 , n21764 );
    not g65 ( n15354 , n2068 );
    not g66 ( n16123 , n25291 );
    and g67 ( n13123 , n8434 , n12016 );
    not g68 ( n25558 , n13660 );
    nor g69 ( n4150 , n4334 , n28870 );
    xnor g70 ( n19853 , n13034 , n21735 );
    not g71 ( n23019 , n19194 );
    or g72 ( n26619 , n4152 , n29872 );
    and g73 ( n18269 , n23672 , n7105 );
    not g74 ( n21711 , n18284 );
    and g75 ( n24768 , n1029 , n26053 );
    or g76 ( n11880 , n21918 , n21771 );
    and g77 ( n16038 , n12937 , n25222 );
    nor g78 ( n2384 , n14573 , n15424 );
    nor g79 ( n2685 , n18274 , n26746 );
    not g80 ( n7611 , n23802 );
    or g81 ( n28908 , n16053 , n26323 );
    not g82 ( n1802 , n5147 );
    and g83 ( n11670 , n4503 , n18077 );
    or g84 ( n20248 , n3641 , n27676 );
    not g85 ( n23504 , n29065 );
    xnor g86 ( n4375 , n1173 , n30789 );
    or g87 ( n5828 , n2359 , n26069 );
    xnor g88 ( n10176 , n21202 , n29309 );
    and g89 ( n18026 , n1536 , n26359 );
    xnor g90 ( n18274 , n18021 , n10975 );
    not g91 ( n11730 , n31115 );
    xnor g92 ( n1483 , n8273 , n16238 );
    or g93 ( n16546 , n12333 , n24032 );
    xnor g94 ( n24520 , n1937 , n9998 );
    nor g95 ( n28330 , n28724 , n30321 );
    not g96 ( n19791 , n5013 );
    not g97 ( n10015 , n27758 );
    xnor g98 ( n1896 , n15227 , n24987 );
    nor g99 ( n26336 , n23510 , n28978 );
    or g100 ( n2945 , n16847 , n11648 );
    and g101 ( n15809 , n8250 , n22260 );
    not g102 ( n3037 , n15987 );
    xnor g103 ( n7125 , n29719 , n22787 );
    and g104 ( n22557 , n17403 , n24146 );
    not g105 ( n21956 , n300 );
    not g106 ( n8037 , n26004 );
    not g107 ( n22301 , n19633 );
    and g108 ( n1614 , n18441 , n11292 );
    xnor g109 ( n10974 , n28867 , n20667 );
    or g110 ( n22616 , n4358 , n28906 );
    xnor g111 ( n17510 , n18641 , n8160 );
    or g112 ( n23363 , n21089 , n11777 );
    not g113 ( n4750 , n3106 );
    and g114 ( n25738 , n25767 , n19718 );
    not g115 ( n4124 , n7999 );
    and g116 ( n21129 , n12898 , n13604 );
    not g117 ( n13336 , n20503 );
    not g118 ( n10383 , n18404 );
    xnor g119 ( n10629 , n4864 , n10515 );
    not g120 ( n7503 , n10439 );
    and g121 ( n6823 , n21848 , n13427 );
    xor g122 ( n1159 , n31365 , n18821 );
    and g123 ( n23617 , n27846 , n12376 );
    not g124 ( n15680 , n10255 );
    nor g125 ( n13960 , n16381 , n6707 );
    not g126 ( n14875 , n26665 );
    or g127 ( n23140 , n30996 , n12682 );
    and g128 ( n6057 , n30127 , n5850 );
    nor g129 ( n11153 , n7209 , n31722 );
    or g130 ( n23907 , n7180 , n11102 );
    xnor g131 ( n13358 , n15046 , n15895 );
    or g132 ( n18932 , n7209 , n7488 );
    not g133 ( n11959 , n6141 );
    xnor g134 ( n10122 , n10842 , n7210 );
    and g135 ( n11510 , n24348 , n5087 );
    or g136 ( n17152 , n17851 , n1006 );
    or g137 ( n7197 , n31140 , n29186 );
    nor g138 ( n30532 , n18133 , n731 );
    or g139 ( n16751 , n10813 , n14017 );
    and g140 ( n15015 , n6549 , n12030 );
    not g141 ( n1746 , n1319 );
    not g142 ( n21274 , n7575 );
    or g143 ( n14326 , n13034 , n29129 );
    not g144 ( n260 , n24442 );
    or g145 ( n29333 , n18179 , n25264 );
    and g146 ( n24576 , n3268 , n28856 );
    or g147 ( n27097 , n30252 , n29781 );
    not g148 ( n14124 , n30411 );
    and g149 ( n11168 , n28071 , n4781 );
    or g150 ( n7271 , n5033 , n11766 );
    xnor g151 ( n4979 , n2627 , n1350 );
    and g152 ( n26314 , n17573 , n5762 );
    xor g153 ( n12464 , n22011 , n7030 );
    and g154 ( n6748 , n9687 , n28677 );
    xor g155 ( n25011 , n26979 , n30640 );
    not g156 ( n19699 , n13244 );
    xnor g157 ( n24160 , n16558 , n25089 );
    or g158 ( n30288 , n24246 , n27135 );
    not g159 ( n24989 , n4978 );
    not g160 ( n15873 , n23115 );
    and g161 ( n14152 , n26704 , n11930 );
    not g162 ( n21446 , n5525 );
    xnor g163 ( n4056 , n5304 , n22567 );
    or g164 ( n8634 , n9876 , n8556 );
    nor g165 ( n15769 , n29080 , n30087 );
    or g166 ( n2132 , n20675 , n17881 );
    xnor g167 ( n24804 , n22812 , n8770 );
    or g168 ( n3114 , n30230 , n997 );
    xnor g169 ( n20927 , n20633 , n11237 );
    nor g170 ( n9981 , n13493 , n27837 );
    and g171 ( n4762 , n19230 , n20725 );
    and g172 ( n11359 , n13258 , n30827 );
    xnor g173 ( n19666 , n18316 , n18030 );
    or g174 ( n24723 , n6969 , n966 );
    or g175 ( n8635 , n2825 , n2225 );
    not g176 ( n17025 , n11177 );
    not g177 ( n29114 , n9241 );
    not g178 ( n3606 , n14235 );
    xnor g179 ( n13181 , n14886 , n18424 );
    not g180 ( n25773 , n9359 );
    not g181 ( n19373 , n2443 );
    and g182 ( n7785 , n591 , n24396 );
    and g183 ( n24659 , n27950 , n17422 );
    and g184 ( n15823 , n29224 , n5685 );
    or g185 ( n22703 , n828 , n3595 );
    and g186 ( n4416 , n13787 , n13053 );
    and g187 ( n29158 , n30587 , n614 );
    nor g188 ( n27813 , n5783 , n19754 );
    xnor g189 ( n12038 , n29775 , n18393 );
    or g190 ( n23264 , n28802 , n29081 );
    or g191 ( n14365 , n460 , n7057 );
    xnor g192 ( n14603 , n23393 , n24242 );
    and g193 ( n5881 , n26202 , n30096 );
    not g194 ( n7423 , n10416 );
    xnor g195 ( n8419 , n14100 , n29615 );
    nor g196 ( n18289 , n30061 , n14618 );
    not g197 ( n30216 , n14888 );
    xnor g198 ( n16414 , n3435 , n6256 );
    xnor g199 ( n7776 , n8199 , n12862 );
    or g200 ( n745 , n25564 , n1804 );
    and g201 ( n20340 , n25992 , n17806 );
    not g202 ( n2690 , n1424 );
    or g203 ( n6441 , n24155 , n30315 );
    not g204 ( n22246 , n7470 );
    not g205 ( n15639 , n5866 );
    not g206 ( n7469 , n17644 );
    not g207 ( n6658 , n10083 );
    and g208 ( n29147 , n25240 , n7008 );
    or g209 ( n10039 , n19300 , n7857 );
    and g210 ( n24269 , n13439 , n10339 );
    not g211 ( n8471 , n21215 );
    xnor g212 ( n24666 , n3421 , n16484 );
    or g213 ( n31760 , n18819 , n22067 );
    xnor g214 ( n10966 , n7667 , n5055 );
    xnor g215 ( n20276 , n16974 , n25666 );
    not g216 ( n11332 , n10238 );
    or g217 ( n12432 , n19398 , n15670 );
    not g218 ( n30428 , n21940 );
    or g219 ( n819 , n7765 , n7933 );
    and g220 ( n22820 , n26223 , n19037 );
    not g221 ( n9933 , n17183 );
    and g222 ( n8734 , n28053 , n3467 );
    not g223 ( n2032 , n12728 );
    xnor g224 ( n29947 , n26315 , n13743 );
    or g225 ( n8829 , n21387 , n10110 );
    or g226 ( n25967 , n2170 , n26830 );
    not g227 ( n15876 , n23101 );
    or g228 ( n24197 , n12348 , n20824 );
    or g229 ( n6671 , n30772 , n16624 );
    not g230 ( n13951 , n18811 );
    and g231 ( n18698 , n16784 , n17823 );
    xnor g232 ( n4799 , n31434 , n25783 );
    or g233 ( n27280 , n13325 , n29637 );
    or g234 ( n5994 , n26078 , n3412 );
    or g235 ( n19271 , n21854 , n7821 );
    not g236 ( n4093 , n25220 );
    nor g237 ( n25534 , n3873 , n346 );
    xor g238 ( n11323 , n3490 , n28405 );
    or g239 ( n8262 , n25069 , n13724 );
    not g240 ( n24471 , n29990 );
    xnor g241 ( n9182 , n11462 , n13604 );
    xnor g242 ( n7502 , n19553 , n22794 );
    nor g243 ( n11486 , n18388 , n30685 );
    not g244 ( n25735 , n12640 );
    not g245 ( n18723 , n29296 );
    and g246 ( n25111 , n4076 , n9692 );
    xnor g247 ( n30961 , n30234 , n2483 );
    or g248 ( n17870 , n1095 , n18550 );
    xnor g249 ( n9781 , n4339 , n29764 );
    and g250 ( n28478 , n4518 , n11221 );
    and g251 ( n31245 , n21348 , n3317 );
    not g252 ( n14994 , n11289 );
    not g253 ( n21038 , n12478 );
    xnor g254 ( n28936 , n10389 , n8865 );
    xnor g255 ( n1361 , n22563 , n4532 );
    or g256 ( n16247 , n26021 , n17070 );
    not g257 ( n7342 , n20305 );
    and g258 ( n22484 , n22160 , n2475 );
    not g259 ( n29484 , n25460 );
    or g260 ( n1689 , n18195 , n15248 );
    not g261 ( n26181 , n20917 );
    nor g262 ( n15367 , n14359 , n17730 );
    nor g263 ( n15645 , n27704 , n14463 );
    nor g264 ( n23601 , n10368 , n20755 );
    xnor g265 ( n924 , n5785 , n13841 );
    not g266 ( n32008 , n3498 );
    and g267 ( n6825 , n5772 , n26918 );
    and g268 ( n10135 , n31430 , n18998 );
    and g269 ( n31345 , n4249 , n25103 );
    nor g270 ( n5799 , n14967 , n7457 );
    and g271 ( n987 , n26520 , n23272 );
    or g272 ( n22621 , n8348 , n25798 );
    or g273 ( n6635 , n14684 , n29263 );
    not g274 ( n11300 , n29435 );
    xnor g275 ( n4959 , n14283 , n23630 );
    not g276 ( n23963 , n4032 );
    or g277 ( n878 , n27331 , n9294 );
    not g278 ( n10271 , n29345 );
    or g279 ( n24447 , n30473 , n17153 );
    and g280 ( n2678 , n4401 , n10415 );
    not g281 ( n14425 , n31098 );
    nor g282 ( n23439 , n19485 , n7772 );
    nor g283 ( n5751 , n23423 , n2357 );
    or g284 ( n28383 , n3488 , n15190 );
    xnor g285 ( n29409 , n7483 , n24223 );
    not g286 ( n5642 , n5271 );
    xnor g287 ( n19270 , n285 , n18259 );
    not g288 ( n21480 , n4172 );
    or g289 ( n12842 , n15606 , n27788 );
    nor g290 ( n17839 , n664 , n17255 );
    not g291 ( n30943 , n13454 );
    or g292 ( n18522 , n16317 , n21413 );
    xnor g293 ( n5854 , n28309 , n18637 );
    and g294 ( n23466 , n30424 , n3255 );
    xnor g295 ( n10142 , n20729 , n5300 );
    or g296 ( n783 , n8905 , n1239 );
    or g297 ( n23376 , n20453 , n8722 );
    not g298 ( n11590 , n31786 );
    or g299 ( n24316 , n16443 , n16429 );
    xnor g300 ( n20084 , n23942 , n1485 );
    and g301 ( n8377 , n21609 , n8493 );
    or g302 ( n27976 , n2225 , n19227 );
    or g303 ( n5950 , n5169 , n4231 );
    xnor g304 ( n25495 , n4823 , n19302 );
    not g305 ( n21544 , n10981 );
    or g306 ( n15344 , n27637 , n546 );
    or g307 ( n12197 , n19524 , n23430 );
    not g308 ( n31845 , n18462 );
    not g309 ( n22714 , n20333 );
    nor g310 ( n21206 , n10681 , n26707 );
    nor g311 ( n30211 , n8111 , n9852 );
    and g312 ( n26521 , n11454 , n7436 );
    and g313 ( n20951 , n11337 , n20016 );
    not g314 ( n10682 , n24255 );
    xnor g315 ( n31568 , n29481 , n25911 );
    not g316 ( n21384 , n31725 );
    and g317 ( n3341 , n16060 , n22445 );
    not g318 ( n20601 , n13975 );
    or g319 ( n11173 , n23892 , n30016 );
    not g320 ( n13790 , n28135 );
    xnor g321 ( n6815 , n9983 , n28988 );
    xnor g322 ( n28121 , n31846 , n19309 );
    and g323 ( n16097 , n11757 , n19413 );
    xnor g324 ( n16610 , n5992 , n7804 );
    or g325 ( n9990 , n3934 , n6976 );
    not g326 ( n23891 , n22804 );
    and g327 ( n15851 , n14164 , n12650 );
    buf g328 ( n6422 , n8356 );
    or g329 ( n22310 , n12871 , n31425 );
    nor g330 ( n20557 , n25436 , n8505 );
    xnor g331 ( n7932 , n15437 , n24743 );
    xnor g332 ( n15572 , n3980 , n16411 );
    xnor g333 ( n24473 , n1243 , n25691 );
    xnor g334 ( n14977 , n23010 , n27570 );
    xnor g335 ( n20848 , n31874 , n8401 );
    or g336 ( n22605 , n8097 , n17590 );
    xnor g337 ( n15592 , n27399 , n20407 );
    xnor g338 ( n16705 , n22130 , n21832 );
    or g339 ( n23478 , n11177 , n19885 );
    or g340 ( n15821 , n27679 , n25802 );
    not g341 ( n4996 , n2060 );
    and g342 ( n8461 , n1928 , n11638 );
    xnor g343 ( n7150 , n4857 , n13105 );
    not g344 ( n3592 , n223 );
    not g345 ( n8436 , n27860 );
    or g346 ( n9922 , n16537 , n14592 );
    and g347 ( n8858 , n16065 , n5647 );
    nor g348 ( n13010 , n20236 , n15142 );
    xnor g349 ( n5794 , n30466 , n22618 );
    not g350 ( n14556 , n24828 );
    xnor g351 ( n22633 , n14218 , n19057 );
    or g352 ( n10950 , n11378 , n9658 );
    or g353 ( n24759 , n18825 , n12672 );
    or g354 ( n12461 , n26677 , n4088 );
    and g355 ( n13426 , n29007 , n9148 );
    not g356 ( n14744 , n14423 );
    xnor g357 ( n23598 , n10936 , n9769 );
    or g358 ( n6908 , n9165 , n907 );
    not g359 ( n22166 , n7389 );
    not g360 ( n8120 , n8042 );
    not g361 ( n25162 , n12821 );
    not g362 ( n3789 , n1823 );
    or g363 ( n25658 , n2025 , n93 );
    and g364 ( n19963 , n30001 , n14234 );
    or g365 ( n7105 , n5963 , n31519 );
    nor g366 ( n13236 , n27089 , n25027 );
    not g367 ( n13761 , n17761 );
    or g368 ( n6219 , n30368 , n4948 );
    xnor g369 ( n4936 , n23875 , n22085 );
    not g370 ( n6698 , n30293 );
    and g371 ( n1799 , n31008 , n24227 );
    or g372 ( n29191 , n15025 , n18828 );
    or g373 ( n16722 , n28863 , n31858 );
    xnor g374 ( n16788 , n352 , n8264 );
    or g375 ( n28295 , n15791 , n10187 );
    or g376 ( n30542 , n16962 , n748 );
    xnor g377 ( n7529 , n19240 , n13271 );
    xnor g378 ( n8434 , n22627 , n22763 );
    xnor g379 ( n26198 , n9284 , n5076 );
    not g380 ( n17209 , n20171 );
    or g381 ( n31351 , n23034 , n20742 );
    xnor g382 ( n12449 , n11140 , n20080 );
    xnor g383 ( n18019 , n1262 , n7227 );
    and g384 ( n2507 , n6227 , n14804 );
    and g385 ( n15054 , n5756 , n17892 );
    not g386 ( n8274 , n29764 );
    or g387 ( n14358 , n15000 , n21602 );
    and g388 ( n29995 , n23812 , n27642 );
    or g389 ( n5624 , n24640 , n18150 );
    not g390 ( n887 , n812 );
    xnor g391 ( n22731 , n6958 , n18622 );
    or g392 ( n23904 , n10440 , n12836 );
    and g393 ( n13996 , n13875 , n25546 );
    nor g394 ( n2698 , n8745 , n23216 );
    not g395 ( n22723 , n16053 );
    not g396 ( n9354 , n4804 );
    or g397 ( n10877 , n678 , n3224 );
    or g398 ( n22063 , n8112 , n23497 );
    or g399 ( n15203 , n24175 , n27995 );
    or g400 ( n6292 , n17571 , n28051 );
    xnor g401 ( n5937 , n15764 , n29538 );
    not g402 ( n2268 , n13688 );
    or g403 ( n10581 , n21173 , n6818 );
    not g404 ( n998 , n454 );
    or g405 ( n24565 , n17873 , n49 );
    and g406 ( n18285 , n13100 , n3381 );
    or g407 ( n1517 , n28254 , n30053 );
    or g408 ( n3751 , n18611 , n14194 );
    not g409 ( n8013 , n6840 );
    xnor g410 ( n21749 , n23807 , n18958 );
    and g411 ( n31720 , n17248 , n23040 );
    not g412 ( n10406 , n22238 );
    not g413 ( n1803 , n4219 );
    xnor g414 ( n16552 , n9742 , n28131 );
    not g415 ( n23897 , n1819 );
    xnor g416 ( n13621 , n26052 , n22675 );
    not g417 ( n20739 , n5652 );
    or g418 ( n3219 , n15583 , n22732 );
    xnor g419 ( n8711 , n13185 , n27974 );
    xnor g420 ( n9949 , n24522 , n20881 );
    and g421 ( n13624 , n31902 , n15203 );
    xor g422 ( n8503 , n27343 , n27688 );
    not g423 ( n21432 , n6253 );
    xnor g424 ( n20514 , n18085 , n6112 );
    and g425 ( n26651 , n21880 , n3086 );
    and g426 ( n7065 , n14932 , n29541 );
    nor g427 ( n29295 , n10028 , n18533 );
    xnor g428 ( n31466 , n2124 , n16643 );
    not g429 ( n10165 , n4423 );
    nor g430 ( n14947 , n5873 , n18389 );
    and g431 ( n13544 , n18573 , n970 );
    or g432 ( n14244 , n22199 , n13337 );
    xnor g433 ( n235 , n25167 , n17917 );
    not g434 ( n1139 , n823 );
    or g435 ( n4035 , n15210 , n30945 );
    and g436 ( n27841 , n28706 , n24912 );
    not g437 ( n20713 , n3626 );
    or g438 ( n21543 , n11885 , n15277 );
    or g439 ( n28651 , n12366 , n21054 );
    and g440 ( n15898 , n12868 , n11006 );
    xnor g441 ( n9610 , n7728 , n7707 );
    not g442 ( n2328 , n19036 );
    not g443 ( n9881 , n3600 );
    xnor g444 ( n17124 , n17368 , n28433 );
    or g445 ( n18406 , n21478 , n18168 );
    not g446 ( n9877 , n31231 );
    or g447 ( n31852 , n6629 , n26267 );
    and g448 ( n21335 , n14115 , n22097 );
    or g449 ( n28506 , n15812 , n2423 );
    xnor g450 ( n24245 , n22405 , n27718 );
    and g451 ( n13499 , n23239 , n30478 );
    not g452 ( n5696 , n28545 );
    or g453 ( n6903 , n8733 , n338 );
    not g454 ( n30486 , n23934 );
    or g455 ( n20331 , n27816 , n25547 );
    and g456 ( n28396 , n26501 , n3532 );
    and g457 ( n14607 , n5980 , n22048 );
    and g458 ( n14686 , n30657 , n10118 );
    not g459 ( n28654 , n29898 );
    nor g460 ( n8682 , n9807 , n22743 );
    or g461 ( n25221 , n3452 , n18154 );
    or g462 ( n22321 , n26025 , n13228 );
    and g463 ( n31804 , n27773 , n6205 );
    not g464 ( n26828 , n9865 );
    or g465 ( n14228 , n27443 , n30826 );
    nor g466 ( n9491 , n10385 , n21719 );
    not g467 ( n21302 , n23773 );
    or g468 ( n9489 , n13903 , n8358 );
    not g469 ( n2508 , n16412 );
    nor g470 ( n14457 , n31481 , n13535 );
    not g471 ( n31185 , n22381 );
    not g472 ( n6419 , n29948 );
    not g473 ( n30939 , n18731 );
    not g474 ( n8164 , n3513 );
    not g475 ( n10439 , n12727 );
    xnor g476 ( n25960 , n26191 , n17910 );
    xnor g477 ( n9350 , n23383 , n30114 );
    or g478 ( n6161 , n24177 , n9504 );
    and g479 ( n22406 , n30858 , n4048 );
    and g480 ( n21732 , n8129 , n30361 );
    not g481 ( n6866 , n24703 );
    xnor g482 ( n3573 , n4444 , n4979 );
    and g483 ( n5351 , n29557 , n17148 );
    or g484 ( n25522 , n5887 , n7292 );
    not g485 ( n14432 , n30002 );
    xnor g486 ( n13984 , n1642 , n24262 );
    nor g487 ( n21752 , n28201 , n2386 );
    not g488 ( n34 , n2018 );
    xor g489 ( n2058 , n21360 , n9709 );
    or g490 ( n10096 , n4756 , n30979 );
    xnor g491 ( n16462 , n19201 , n20214 );
    nor g492 ( n2280 , n30238 , n26534 );
    nor g493 ( n24297 , n20881 , n15559 );
    nor g494 ( n13255 , n19189 , n19444 );
    and g495 ( n29496 , n7685 , n18521 );
    not g496 ( n26545 , n11931 );
    not g497 ( n15708 , n3416 );
    not g498 ( n11975 , n2405 );
    not g499 ( n16598 , n11658 );
    nor g500 ( n20534 , n27534 , n21443 );
    not g501 ( n9151 , n13561 );
    or g502 ( n10948 , n20256 , n30745 );
    not g503 ( n27239 , n18667 );
    not g504 ( n7052 , n15857 );
    buf g505 ( n25579 , n29393 );
    and g506 ( n24405 , n2746 , n24798 );
    or g507 ( n522 , n20409 , n23535 );
    xnor g508 ( n30815 , n16062 , n23502 );
    or g509 ( n11176 , n27262 , n30654 );
    not g510 ( n21110 , n17478 );
    or g511 ( n3181 , n16326 , n27397 );
    or g512 ( n8916 , n4551 , n21232 );
    or g513 ( n30854 , n30184 , n31165 );
    xnor g514 ( n8354 , n9550 , n1781 );
    not g515 ( n29197 , n29053 );
    and g516 ( n14674 , n3561 , n29913 );
    xnor g517 ( n24781 , n27546 , n19592 );
    not g518 ( n31010 , n24275 );
    and g519 ( n6562 , n2284 , n20094 );
    not g520 ( n22850 , n24481 );
    xnor g521 ( n8046 , n28307 , n7992 );
    not g522 ( n27722 , n20616 );
    and g523 ( n10920 , n4407 , n4171 );
    or g524 ( n10811 , n23188 , n14439 );
    xnor g525 ( n7864 , n31067 , n5685 );
    and g526 ( n17097 , n10948 , n10976 );
    or g527 ( n3625 , n21055 , n184 );
    and g528 ( n31371 , n29747 , n23138 );
    nor g529 ( n1690 , n28189 , n6825 );
    or g530 ( n29468 , n2770 , n6050 );
    or g531 ( n8761 , n3577 , n17578 );
    or g532 ( n1184 , n28699 , n20938 );
    or g533 ( n2402 , n23018 , n31879 );
    or g534 ( n24461 , n9343 , n6745 );
    or g535 ( n334 , n28646 , n24080 );
    nor g536 ( n22538 , n20390 , n28829 );
    and g537 ( n14428 , n3900 , n9140 );
    xnor g538 ( n29398 , n3450 , n11056 );
    nor g539 ( n14535 , n1285 , n30593 );
    or g540 ( n3538 , n11354 , n15934 );
    nor g541 ( n20128 , n13632 , n19791 );
    not g542 ( n27967 , n16080 );
    not g543 ( n17682 , n26237 );
    not g544 ( n18431 , n30696 );
    not g545 ( n24762 , n5781 );
    nor g546 ( n27028 , n8364 , n29839 );
    xnor g547 ( n6089 , n11593 , n21971 );
    xnor g548 ( n14013 , n25942 , n18369 );
    or g549 ( n17392 , n26535 , n30415 );
    nor g550 ( n30092 , n17557 , n13634 );
    not g551 ( n26659 , n6419 );
    not g552 ( n914 , n7482 );
    xnor g553 ( n6937 , n31876 , n21008 );
    or g554 ( n12376 , n16942 , n11918 );
    xnor g555 ( n13424 , n30074 , n14817 );
    not g556 ( n11188 , n4760 );
    xnor g557 ( n20871 , n28204 , n17843 );
    xnor g558 ( n14984 , n3014 , n124 );
    or g559 ( n8755 , n124 , n15027 );
    and g560 ( n12796 , n25601 , n7274 );
    not g561 ( n26179 , n26403 );
    or g562 ( n18991 , n13578 , n4546 );
    xnor g563 ( n404 , n31410 , n26474 );
    nor g564 ( n30860 , n22555 , n16004 );
    xnor g565 ( n982 , n25210 , n25915 );
    nor g566 ( n7754 , n21261 , n21963 );
    or g567 ( n7477 , n26018 , n11582 );
    or g568 ( n3227 , n9875 , n2503 );
    xnor g569 ( n25935 , n6670 , n12967 );
    xnor g570 ( n29988 , n26495 , n29176 );
    xnor g571 ( n14079 , n19564 , n2799 );
    nor g572 ( n5852 , n27948 , n4771 );
    nor g573 ( n9133 , n3505 , n3710 );
    not g574 ( n13518 , n20144 );
    or g575 ( n12372 , n31094 , n114 );
    nor g576 ( n7714 , n8867 , n26696 );
    or g577 ( n26881 , n2826 , n1211 );
    not g578 ( n18948 , n11833 );
    or g579 ( n9009 , n21626 , n17256 );
    or g580 ( n17576 , n2843 , n16580 );
    nor g581 ( n26240 , n22349 , n13417 );
    xnor g582 ( n19302 , n11427 , n21161 );
    xnor g583 ( n12308 , n14785 , n6541 );
    or g584 ( n14530 , n30020 , n5326 );
    not g585 ( n8550 , n19717 );
    or g586 ( n3035 , n12251 , n2301 );
    nor g587 ( n17869 , n18907 , n1995 );
    xnor g588 ( n778 , n13814 , n20587 );
    xnor g589 ( n19173 , n12625 , n21185 );
    and g590 ( n26563 , n16666 , n12621 );
    not g591 ( n29656 , n4374 );
    xnor g592 ( n13781 , n13716 , n8370 );
    or g593 ( n18588 , n24225 , n13791 );
    xnor g594 ( n26669 , n22229 , n2828 );
    or g595 ( n2161 , n10433 , n2842 );
    nor g596 ( n29911 , n7547 , n10524 );
    xnor g597 ( n13149 , n16777 , n11948 );
    xnor g598 ( n10325 , n30184 , n12162 );
    or g599 ( n253 , n12857 , n7338 );
    or g600 ( n5878 , n8473 , n19293 );
    nor g601 ( n7836 , n16441 , n1414 );
    and g602 ( n21202 , n9841 , n15330 );
    xnor g603 ( n16852 , n15008 , n13256 );
    not g604 ( n7369 , n31323 );
    or g605 ( n3721 , n2065 , n26740 );
    not g606 ( n29431 , n3540 );
    nor g607 ( n2206 , n1995 , n24920 );
    or g608 ( n27516 , n20309 , n8182 );
    not g609 ( n1229 , n18871 );
    not g610 ( n30401 , n28815 );
    nor g611 ( n5568 , n6936 , n28809 );
    not g612 ( n29960 , n23398 );
    xnor g613 ( n29816 , n12604 , n2178 );
    and g614 ( n29820 , n5868 , n19274 );
    and g615 ( n29430 , n7348 , n11166 );
    not g616 ( n3427 , n11361 );
    not g617 ( n16970 , n3198 );
    and g618 ( n19740 , n7603 , n20276 );
    not g619 ( n14841 , n3867 );
    nor g620 ( n25180 , n18378 , n386 );
    not g621 ( n10150 , n19091 );
    and g622 ( n23196 , n31983 , n17991 );
    nor g623 ( n25556 , n3043 , n19029 );
    or g624 ( n31208 , n26715 , n308 );
    xnor g625 ( n30188 , n16738 , n22642 );
    not g626 ( n23201 , n5803 );
    or g627 ( n22526 , n7434 , n15142 );
    or g628 ( n2304 , n2024 , n30865 );
    nor g629 ( n17014 , n21032 , n27892 );
    and g630 ( n28992 , n25862 , n8030 );
    xnor g631 ( n24905 , n12039 , n8130 );
    and g632 ( n29260 , n3601 , n2593 );
    or g633 ( n14440 , n3081 , n6245 );
    not g634 ( n26219 , n28742 );
    and g635 ( n7829 , n543 , n13709 );
    xnor g636 ( n10593 , n6159 , n14896 );
    or g637 ( n4437 , n10276 , n19684 );
    not g638 ( n27401 , n20914 );
    or g639 ( n3623 , n1943 , n8766 );
    xnor g640 ( n22224 , n15536 , n6777 );
    and g641 ( n8985 , n12573 , n23097 );
    xor g642 ( n26807 , n12556 , n2550 );
    not g643 ( n31249 , n417 );
    not g644 ( n724 , n29380 );
    or g645 ( n13085 , n9757 , n5459 );
    or g646 ( n3074 , n16712 , n19626 );
    xnor g647 ( n8532 , n23852 , n28562 );
    and g648 ( n7649 , n3760 , n15021 );
    xnor g649 ( n29547 , n5859 , n3365 );
    or g650 ( n17137 , n3896 , n14211 );
    not g651 ( n15525 , n30141 );
    or g652 ( n11077 , n20000 , n7774 );
    and g653 ( n7416 , n6219 , n7430 );
    or g654 ( n13027 , n4408 , n29645 );
    or g655 ( n10547 , n10322 , n4102 );
    or g656 ( n3671 , n29510 , n28003 );
    xnor g657 ( n11331 , n3345 , n16516 );
    and g658 ( n19938 , n27122 , n30593 );
    nor g659 ( n29020 , n2719 , n12910 );
    and g660 ( n29235 , n25658 , n2104 );
    or g661 ( n12549 , n22736 , n14449 );
    and g662 ( n19927 , n19863 , n13550 );
    and g663 ( n24421 , n3738 , n697 );
    or g664 ( n4937 , n13487 , n8012 );
    nor g665 ( n2645 , n30409 , n10154 );
    not g666 ( n25253 , n30642 );
    or g667 ( n5522 , n2780 , n2036 );
    xnor g668 ( n16328 , n14855 , n359 );
    xnor g669 ( n21098 , n24236 , n22845 );
    and g670 ( n3402 , n5872 , n8591 );
    not g671 ( n28979 , n2150 );
    nor g672 ( n14782 , n21064 , n20057 );
    xnor g673 ( n3956 , n30194 , n10118 );
    buf g674 ( n1331 , n121 );
    not g675 ( n16218 , n14004 );
    not g676 ( n30687 , n12130 );
    not g677 ( n21896 , n22306 );
    or g678 ( n15768 , n1195 , n26005 );
    buf g679 ( n20412 , n26186 );
    nor g680 ( n27980 , n14324 , n10861 );
    nor g681 ( n31558 , n26691 , n4969 );
    and g682 ( n9664 , n9008 , n5251 );
    or g683 ( n29749 , n16362 , n30144 );
    not g684 ( n21685 , n449 );
    or g685 ( n20277 , n28259 , n13574 );
    not g686 ( n25298 , n16171 );
    and g687 ( n28232 , n13567 , n2737 );
    and g688 ( n1622 , n745 , n22729 );
    not g689 ( n5574 , n25162 );
    xnor g690 ( n7148 , n25475 , n5968 );
    not g691 ( n14751 , n24377 );
    xnor g692 ( n20768 , n26818 , n535 );
    or g693 ( n10372 , n2656 , n9533 );
    not g694 ( n18000 , n8264 );
    or g695 ( n18872 , n23327 , n17675 );
    buf g696 ( n30321 , n16077 );
    not g697 ( n8308 , n31783 );
    xnor g698 ( n32 , n9513 , n15006 );
    not g699 ( n485 , n15689 );
    nor g700 ( n15441 , n11517 , n10454 );
    or g701 ( n32022 , n22131 , n27107 );
    or g702 ( n20654 , n12968 , n976 );
    xnor g703 ( n13498 , n215 , n20905 );
    not g704 ( n31431 , n19861 );
    or g705 ( n16658 , n25008 , n29628 );
    xnor g706 ( n5001 , n23015 , n16370 );
    or g707 ( n247 , n16424 , n30259 );
    nor g708 ( n533 , n13575 , n11857 );
    not g709 ( n9270 , n29741 );
    not g710 ( n16483 , n20786 );
    or g711 ( n17534 , n9910 , n26345 );
    and g712 ( n3146 , n22797 , n11783 );
    or g713 ( n12203 , n27275 , n18242 );
    xnor g714 ( n23536 , n25345 , n28572 );
    not g715 ( n537 , n1283 );
    xnor g716 ( n16484 , n22246 , n22355 );
    buf g717 ( n6882 , n6883 );
    not g718 ( n17380 , n7010 );
    not g719 ( n21197 , n11563 );
    and g720 ( n31799 , n4633 , n3969 );
    not g721 ( n1100 , n28081 );
    or g722 ( n40 , n5826 , n29616 );
    xnor g723 ( n11935 , n12670 , n21315 );
    not g724 ( n20078 , n5160 );
    not g725 ( n17653 , n26290 );
    not g726 ( n13934 , n6082 );
    xnor g727 ( n27678 , n25399 , n31204 );
    not g728 ( n17243 , n8613 );
    not g729 ( n4904 , n10398 );
    or g730 ( n25363 , n17143 , n5465 );
    not g731 ( n31743 , n6639 );
    nor g732 ( n31147 , n13604 , n5456 );
    or g733 ( n24227 , n7147 , n20105 );
    or g734 ( n809 , n28203 , n26005 );
    xnor g735 ( n18131 , n29297 , n12806 );
    not g736 ( n6243 , n17109 );
    and g737 ( n13497 , n11765 , n20561 );
    and g738 ( n15736 , n18029 , n626 );
    not g739 ( n19999 , n891 );
    and g740 ( n14824 , n15290 , n20821 );
    or g741 ( n26936 , n18875 , n18364 );
    nor g742 ( n3051 , n17068 , n6349 );
    nor g743 ( n13274 , n18669 , n1770 );
    nor g744 ( n6132 , n8986 , n5313 );
    and g745 ( n13449 , n28892 , n27154 );
    not g746 ( n13992 , n18966 );
    and g747 ( n3550 , n1909 , n26252 );
    or g748 ( n1750 , n12795 , n3908 );
    not g749 ( n1931 , n29168 );
    not g750 ( n23127 , n13768 );
    and g751 ( n26393 , n28286 , n28326 );
    xnor g752 ( n10990 , n25602 , n12508 );
    xnor g753 ( n21625 , n14809 , n1883 );
    not g754 ( n19332 , n3238 );
    xnor g755 ( n20169 , n3967 , n30201 );
    nor g756 ( n3663 , n3432 , n1078 );
    xnor g757 ( n4972 , n24184 , n29059 );
    and g758 ( n25231 , n1757 , n16704 );
    and g759 ( n17578 , n23860 , n8744 );
    nor g760 ( n4006 , n23043 , n15807 );
    not g761 ( n5936 , n19248 );
    xnor g762 ( n4419 , n19520 , n29045 );
    or g763 ( n6994 , n19348 , n5261 );
    or g764 ( n31716 , n6874 , n6596 );
    and g765 ( n30051 , n26724 , n10008 );
    or g766 ( n2812 , n25551 , n29196 );
    not g767 ( n25061 , n31591 );
    and g768 ( n7415 , n25662 , n2276 );
    xnor g769 ( n23542 , n17598 , n1579 );
    not g770 ( n14400 , n1191 );
    buf g771 ( n6745 , n28378 );
    and g772 ( n21152 , n1607 , n4211 );
    and g773 ( n19081 , n7495 , n20155 );
    nor g774 ( n10645 , n20728 , n4929 );
    or g775 ( n11961 , n19764 , n24157 );
    or g776 ( n22908 , n24124 , n426 );
    not g777 ( n22336 , n5011 );
    not g778 ( n27512 , n3486 );
    xnor g779 ( n7151 , n17690 , n18620 );
    nor g780 ( n10333 , n27077 , n17884 );
    not g781 ( n9301 , n22994 );
    xnor g782 ( n10706 , n14510 , n22434 );
    and g783 ( n6907 , n28651 , n11542 );
    xnor g784 ( n15417 , n12301 , n21475 );
    xnor g785 ( n4645 , n19268 , n17917 );
    not g786 ( n12764 , n3565 );
    xnor g787 ( n27676 , n4486 , n17251 );
    nor g788 ( n3987 , n626 , n24621 );
    or g789 ( n26478 , n23427 , n4475 );
    and g790 ( n3258 , n28184 , n10478 );
    or g791 ( n20520 , n18785 , n17056 );
    xnor g792 ( n6270 , n25899 , n3962 );
    xnor g793 ( n3820 , n29380 , n12398 );
    not g794 ( n7718 , n28633 );
    or g795 ( n16020 , n21636 , n10653 );
    and g796 ( n4462 , n11639 , n13685 );
    xor g797 ( n8622 , n9725 , n3268 );
    nor g798 ( n16012 , n26324 , n29881 );
    xnor g799 ( n14470 , n30936 , n20736 );
    or g800 ( n12611 , n1568 , n12402 );
    not g801 ( n27844 , n15152 );
    not g802 ( n19935 , n23195 );
    and g803 ( n4256 , n28501 , n8873 );
    or g804 ( n4903 , n24975 , n26581 );
    xnor g805 ( n6946 , n9149 , n1411 );
    and g806 ( n28183 , n12248 , n30986 );
    not g807 ( n7859 , n28417 );
    or g808 ( n22839 , n19498 , n3674 );
    and g809 ( n29964 , n22383 , n6171 );
    xnor g810 ( n25700 , n8321 , n7209 );
    or g811 ( n9050 , n2528 , n24225 );
    and g812 ( n7419 , n3958 , n13750 );
    and g813 ( n6229 , n6064 , n12635 );
    nor g814 ( n28401 , n29878 , n7560 );
    not g815 ( n25987 , n13391 );
    not g816 ( n26066 , n4836 );
    and g817 ( n15732 , n3464 , n13737 );
    xnor g818 ( n21885 , n12569 , n27741 );
    not g819 ( n29525 , n1724 );
    or g820 ( n23599 , n9505 , n25826 );
    xnor g821 ( n31665 , n25237 , n25838 );
    and g822 ( n5552 , n380 , n9947 );
    xnor g823 ( n22796 , n15039 , n5559 );
    xnor g824 ( n21942 , n17330 , n1635 );
    xnor g825 ( n29804 , n19837 , n8798 );
    and g826 ( n14976 , n5819 , n3214 );
    not g827 ( n12400 , n9575 );
    not g828 ( n17531 , n4412 );
    or g829 ( n16482 , n23400 , n9650 );
    not g830 ( n27826 , n6863 );
    not g831 ( n658 , n21358 );
    nor g832 ( n19554 , n14434 , n2589 );
    not g833 ( n11889 , n12385 );
    or g834 ( n15974 , n29851 , n1678 );
    xnor g835 ( n31127 , n28522 , n10817 );
    or g836 ( n7098 , n1615 , n3341 );
    or g837 ( n19609 , n18165 , n20150 );
    xnor g838 ( n15591 , n13904 , n1144 );
    xnor g839 ( n30391 , n31750 , n20144 );
    or g840 ( n29917 , n12916 , n2585 );
    or g841 ( n562 , n9870 , n15028 );
    and g842 ( n20103 , n27614 , n2448 );
    and g843 ( n2600 , n7185 , n11183 );
    not g844 ( n27994 , n14434 );
    not g845 ( n30106 , n5027 );
    or g846 ( n24955 , n10688 , n21204 );
    or g847 ( n14265 , n19711 , n2200 );
    xnor g848 ( n13520 , n11458 , n26598 );
    xor g849 ( n13677 , n22605 , n862 );
    or g850 ( n30682 , n18132 , n6951 );
    xnor g851 ( n21307 , n27999 , n12974 );
    xnor g852 ( n22813 , n27651 , n25365 );
    nor g853 ( n23795 , n3432 , n5281 );
    not g854 ( n1953 , n7890 );
    or g855 ( n31274 , n19326 , n4827 );
    or g856 ( n9811 , n22628 , n741 );
    or g857 ( n28711 , n17689 , n21532 );
    not g858 ( n3983 , n12760 );
    xor g859 ( n9435 , n30621 , n25538 );
    not g860 ( n13613 , n24086 );
    xnor g861 ( n20766 , n31361 , n13725 );
    or g862 ( n9055 , n2760 , n31195 );
    xnor g863 ( n20455 , n29249 , n20799 );
    xnor g864 ( n16178 , n31060 , n22233 );
    and g865 ( n14341 , n25554 , n29359 );
    not g866 ( n26165 , n23614 );
    not g867 ( n5310 , n20877 );
    or g868 ( n3525 , n26988 , n11458 );
    not g869 ( n17772 , n21670 );
    or g870 ( n14893 , n31241 , n28043 );
    or g871 ( n26113 , n18705 , n10708 );
    or g872 ( n12219 , n28342 , n4381 );
    and g873 ( n3273 , n29333 , n9278 );
    or g874 ( n9093 , n18687 , n30859 );
    xnor g875 ( n29416 , n23809 , n21642 );
    xnor g876 ( n19306 , n21597 , n6957 );
    and g877 ( n20817 , n30413 , n1664 );
    or g878 ( n782 , n27239 , n18216 );
    or g879 ( n6294 , n1022 , n11987 );
    xnor g880 ( n7162 , n19813 , n15869 );
    and g881 ( n27778 , n18264 , n14690 );
    not g882 ( n12912 , n1177 );
    not g883 ( n26804 , n10364 );
    not g884 ( n11286 , n4848 );
    nor g885 ( n31769 , n30201 , n28453 );
    or g886 ( n15473 , n30936 , n20736 );
    xnor g887 ( n31224 , n5034 , n15922 );
    nor g888 ( n18957 , n6171 , n18561 );
    not g889 ( n13817 , n2920 );
    not g890 ( n8486 , n14641 );
    xor g891 ( n15094 , n18694 , n27391 );
    not g892 ( n1412 , n22041 );
    or g893 ( n2623 , n26473 , n2454 );
    xnor g894 ( n5453 , n20175 , n27126 );
    or g895 ( n23917 , n21261 , n22867 );
    not g896 ( n31520 , n31218 );
    not g897 ( n2759 , n21369 );
    and g898 ( n3761 , n12950 , n6079 );
    and g899 ( n4478 , n18644 , n21245 );
    or g900 ( n16063 , n31458 , n11919 );
    xnor g901 ( n13695 , n18395 , n28445 );
    not g902 ( n18913 , n5274 );
    xnor g903 ( n30506 , n28417 , n13137 );
    or g904 ( n17520 , n28081 , n24893 );
    xnor g905 ( n6961 , n24630 , n11736 );
    or g906 ( n25108 , n14959 , n424 );
    xnor g907 ( n23476 , n5598 , n7755 );
    nor g908 ( n1051 , n20611 , n5435 );
    or g909 ( n5507 , n10051 , n10588 );
    and g910 ( n9753 , n25607 , n31903 );
    or g911 ( n10833 , n15843 , n17350 );
    and g912 ( n30881 , n9754 , n18776 );
    nor g913 ( n12174 , n31917 , n31561 );
    xnor g914 ( n2347 , n3219 , n21370 );
    or g915 ( n28996 , n23676 , n10768 );
    xnor g916 ( n15746 , n3259 , n19255 );
    not g917 ( n17007 , n21166 );
    or g918 ( n30718 , n10494 , n4244 );
    xnor g919 ( n20937 , n29982 , n11716 );
    xnor g920 ( n7288 , n26892 , n25624 );
    not g921 ( n28089 , n12478 );
    and g922 ( n24707 , n29653 , n27171 );
    not g923 ( n20154 , n26456 );
    xnor g924 ( n5247 , n23449 , n28020 );
    and g925 ( n20787 , n7817 , n5009 );
    not g926 ( n17963 , n1800 );
    or g927 ( n2839 , n21306 , n2343 );
    or g928 ( n25034 , n31288 , n29368 );
    xnor g929 ( n12571 , n24409 , n12426 );
    not g930 ( n23058 , n6347 );
    not g931 ( n16843 , n20595 );
    not g932 ( n13167 , n16785 );
    xnor g933 ( n26707 , n9038 , n21796 );
    not g934 ( n31560 , n1298 );
    and g935 ( n22519 , n28536 , n24737 );
    nor g936 ( n22552 , n16311 , n2080 );
    not g937 ( n10585 , n10992 );
    and g938 ( n20830 , n24112 , n24101 );
    nor g939 ( n11228 , n2674 , n24725 );
    xnor g940 ( n5076 , n6249 , n8834 );
    xnor g941 ( n8698 , n4180 , n2195 );
    or g942 ( n8793 , n20282 , n3329 );
    and g943 ( n24249 , n28361 , n16027 );
    nor g944 ( n27780 , n19092 , n3184 );
    not g945 ( n6012 , n28262 );
    xnor g946 ( n4920 , n17626 , n3194 );
    and g947 ( n8872 , n29536 , n3518 );
    and g948 ( n15627 , n861 , n20247 );
    xor g949 ( n2885 , n3316 , n25133 );
    or g950 ( n24250 , n14588 , n30395 );
    or g951 ( n6846 , n23493 , n10697 );
    nor g952 ( n7586 , n16860 , n7258 );
    not g953 ( n6415 , n5137 );
    not g954 ( n17754 , n12962 );
    xnor g955 ( n31319 , n20453 , n11886 );
    not g956 ( n1127 , n11307 );
    or g957 ( n11750 , n18170 , n23528 );
    nor g958 ( n20770 , n26254 , n19982 );
    and g959 ( n16419 , n26050 , n29425 );
    not g960 ( n9529 , n4795 );
    xnor g961 ( n6794 , n3442 , n11521 );
    and g962 ( n18458 , n23862 , n20182 );
    xor g963 ( n14178 , n8269 , n3863 );
    not g964 ( n8967 , n21401 );
    and g965 ( n16207 , n6161 , n18299 );
    not g966 ( n7488 , n27453 );
    or g967 ( n7255 , n10453 , n6796 );
    xnor g968 ( n16485 , n4074 , n1752 );
    or g969 ( n6704 , n10386 , n11015 );
    or g970 ( n6537 , n31715 , n8198 );
    or g971 ( n21744 , n9607 , n25355 );
    xnor g972 ( n1932 , n14935 , n10929 );
    nor g973 ( n27039 , n3269 , n10696 );
    or g974 ( n1215 , n30092 , n28196 );
    xnor g975 ( n17589 , n4791 , n31513 );
    and g976 ( n25625 , n1865 , n1331 );
    and g977 ( n14606 , n19147 , n4984 );
    nor g978 ( n18545 , n15948 , n17888 );
    or g979 ( n3236 , n15317 , n26521 );
    or g980 ( n5605 , n23634 , n17774 );
    not g981 ( n1166 , n15387 );
    and g982 ( n5977 , n336 , n4826 );
    xnor g983 ( n7077 , n20498 , n22223 );
    xnor g984 ( n5381 , n28549 , n26605 );
    xnor g985 ( n3803 , n17365 , n13887 );
    or g986 ( n19389 , n22393 , n13346 );
    nor g987 ( n8100 , n25506 , n20780 );
    or g988 ( n26522 , n17682 , n24584 );
    or g989 ( n18188 , n16989 , n4566 );
    xnor g990 ( n9190 , n20280 , n17374 );
    and g991 ( n11681 , n30123 , n3301 );
    xnor g992 ( n3101 , n3200 , n10282 );
    not g993 ( n16256 , n863 );
    not g994 ( n15954 , n12266 );
    or g995 ( n22672 , n15706 , n5396 );
    xnor g996 ( n14135 , n8926 , n26599 );
    and g997 ( n19812 , n9329 , n20478 );
    and g998 ( n18436 , n5534 , n388 );
    xnor g999 ( n5649 , n12304 , n25781 );
    xnor g1000 ( n13944 , n27762 , n1844 );
    or g1001 ( n12304 , n5620 , n11000 );
    and g1002 ( n16286 , n23916 , n21526 );
    xnor g1003 ( n6504 , n6941 , n4764 );
    xnor g1004 ( n18622 , n15085 , n14777 );
    not g1005 ( n10134 , n11763 );
    nor g1006 ( n30880 , n8605 , n1825 );
    not g1007 ( n10600 , n22855 );
    not g1008 ( n10430 , n30245 );
    and g1009 ( n23695 , n1948 , n23254 );
    not g1010 ( n8783 , n27885 );
    or g1011 ( n4855 , n2704 , n25194 );
    nor g1012 ( n5627 , n1021 , n15354 );
    not g1013 ( n20341 , n23095 );
    xnor g1014 ( n9323 , n17762 , n3440 );
    nor g1015 ( n11823 , n20810 , n9416 );
    xnor g1016 ( n13598 , n26562 , n5514 );
    xnor g1017 ( n31069 , n6194 , n31027 );
    and g1018 ( n6530 , n1706 , n9982 );
    xnor g1019 ( n14173 , n23050 , n3939 );
    xnor g1020 ( n4861 , n11415 , n1518 );
    not g1021 ( n13268 , n13519 );
    and g1022 ( n3708 , n6182 , n18606 );
    not g1023 ( n4466 , n4735 );
    nor g1024 ( n14431 , n18753 , n21609 );
    nor g1025 ( n16840 , n2542 , n19364 );
    not g1026 ( n1294 , n6726 );
    or g1027 ( n12575 , n17813 , n6264 );
    or g1028 ( n21920 , n11894 , n9146 );
    xnor g1029 ( n2567 , n10094 , n11363 );
    or g1030 ( n23225 , n26328 , n26213 );
    xnor g1031 ( n8983 , n2216 , n11974 );
    and g1032 ( n4674 , n17529 , n17816 );
    xnor g1033 ( n2109 , n24192 , n8662 );
    not g1034 ( n29840 , n5612 );
    and g1035 ( n12331 , n22810 , n5819 );
    not g1036 ( n16363 , n1527 );
    xnor g1037 ( n27439 , n7946 , n26541 );
    xor g1038 ( n13118 , n18659 , n7905 );
    xnor g1039 ( n24674 , n18697 , n20325 );
    nor g1040 ( n10739 , n6888 , n20940 );
    xnor g1041 ( n14140 , n5191 , n8074 );
    not g1042 ( n22937 , n17004 );
    xnor g1043 ( n9820 , n268 , n13748 );
    or g1044 ( n26147 , n318 , n12370 );
    not g1045 ( n18798 , n24819 );
    xnor g1046 ( n10461 , n14739 , n13444 );
    xnor g1047 ( n1432 , n27194 , n28830 );
    and g1048 ( n9683 , n10801 , n24137 );
    and g1049 ( n20743 , n2076 , n11348 );
    xnor g1050 ( n17829 , n26722 , n2433 );
    not g1051 ( n19386 , n27925 );
    not g1052 ( n22418 , n22264 );
    and g1053 ( n29534 , n8728 , n16618 );
    not g1054 ( n13254 , n25512 );
    or g1055 ( n14229 , n2286 , n13422 );
    not g1056 ( n15789 , n9378 );
    xnor g1057 ( n12486 , n18523 , n28796 );
    not g1058 ( n20339 , n31757 );
    or g1059 ( n2671 , n26596 , n31174 );
    nor g1060 ( n2411 , n3225 , n5715 );
    not g1061 ( n5819 , n22675 );
    and g1062 ( n8103 , n31564 , n19242 );
    xnor g1063 ( n17731 , n16075 , n22922 );
    xnor g1064 ( n27029 , n8418 , n6046 );
    nor g1065 ( n24319 , n14040 , n561 );
    xor g1066 ( n3720 , n1151 , n21664 );
    not g1067 ( n14834 , n25338 );
    not g1068 ( n18429 , n17990 );
    not g1069 ( n5277 , n12123 );
    or g1070 ( n9651 , n6560 , n22525 );
    not g1071 ( n9412 , n17313 );
    not g1072 ( n4059 , n6401 );
    not g1073 ( n17656 , n17537 );
    or g1074 ( n30379 , n16516 , n8807 );
    not g1075 ( n14612 , n9873 );
    not g1076 ( n21562 , n3569 );
    or g1077 ( n7119 , n9167 , n29313 );
    xnor g1078 ( n23748 , n427 , n5194 );
    or g1079 ( n14158 , n21201 , n16913 );
    and g1080 ( n28793 , n5950 , n2484 );
    xnor g1081 ( n26346 , n22391 , n30803 );
    xnor g1082 ( n31373 , n26475 , n17540 );
    not g1083 ( n12690 , n8726 );
    not g1084 ( n26173 , n4002 );
    not g1085 ( n12706 , n24440 );
    nor g1086 ( n18500 , n6553 , n14517 );
    xnor g1087 ( n18514 , n26428 , n562 );
    or g1088 ( n27852 , n4272 , n14502 );
    xnor g1089 ( n8085 , n31463 , n66 );
    xnor g1090 ( n22802 , n8857 , n24794 );
    nor g1091 ( n13076 , n19728 , n7901 );
    and g1092 ( n18646 , n3841 , n29062 );
    xnor g1093 ( n25679 , n22424 , n17464 );
    not g1094 ( n10890 , n29153 );
    or g1095 ( n14143 , n17911 , n27700 );
    or g1096 ( n22821 , n2616 , n14339 );
    or g1097 ( n22661 , n18061 , n23803 );
    or g1098 ( n21887 , n13180 , n3218 );
    not g1099 ( n25447 , n29188 );
    nor g1100 ( n22750 , n2798 , n17499 );
    not g1101 ( n17819 , n441 );
    not g1102 ( n26254 , n5792 );
    xnor g1103 ( n13205 , n18895 , n6534 );
    and g1104 ( n26736 , n28199 , n21611 );
    xnor g1105 ( n27541 , n15438 , n6641 );
    xnor g1106 ( n19960 , n24273 , n9775 );
    or g1107 ( n8799 , n11670 , n20323 );
    or g1108 ( n18256 , n12487 , n2442 );
    not g1109 ( n15305 , n30228 );
    xnor g1110 ( n23922 , n2771 , n25740 );
    and g1111 ( n20044 , n7814 , n21737 );
    xnor g1112 ( n2323 , n20399 , n1951 );
    nor g1113 ( n24013 , n11253 , n30374 );
    not g1114 ( n31152 , n28243 );
    xor g1115 ( n2410 , n4255 , n9663 );
    or g1116 ( n9143 , n27145 , n5619 );
    not g1117 ( n17924 , n26826 );
    xnor g1118 ( n3152 , n1750 , n24050 );
    xnor g1119 ( n11891 , n13383 , n23965 );
    nor g1120 ( n6314 , n12244 , n28235 );
    nor g1121 ( n20650 , n4257 , n6374 );
    nor g1122 ( n20659 , n17413 , n29794 );
    xnor g1123 ( n11761 , n362 , n24241 );
    not g1124 ( n9071 , n23692 );
    not g1125 ( n26769 , n11905 );
    or g1126 ( n19997 , n17849 , n26973 );
    not g1127 ( n23995 , n757 );
    and g1128 ( n24499 , n22201 , n19565 );
    xnor g1129 ( n15710 , n28442 , n1251 );
    or g1130 ( n18750 , n13949 , n14237 );
    xnor g1131 ( n15500 , n18350 , n30245 );
    not g1132 ( n13061 , n16319 );
    or g1133 ( n23847 , n18649 , n15958 );
    xnor g1134 ( n571 , n563 , n255 );
    not g1135 ( n4791 , n17270 );
    not g1136 ( n5304 , n372 );
    not g1137 ( n13295 , n4426 );
    not g1138 ( n19942 , n138 );
    and g1139 ( n5598 , n30710 , n5684 );
    or g1140 ( n17290 , n24304 , n8187 );
    xnor g1141 ( n2663 , n20236 , n12668 );
    not g1142 ( n31781 , n21757 );
    xnor g1143 ( n31055 , n12152 , n31811 );
    or g1144 ( n7002 , n19167 , n11851 );
    xnor g1145 ( n31904 , n25612 , n14635 );
    xor g1146 ( n24490 , n16769 , n12310 );
    nor g1147 ( n2706 , n25104 , n26176 );
    not g1148 ( n4570 , n22124 );
    or g1149 ( n22356 , n4298 , n14373 );
    not g1150 ( n14708 , n12346 );
    not g1151 ( n11302 , n8584 );
    and g1152 ( n19623 , n11029 , n4321 );
    or g1153 ( n17401 , n13845 , n8928 );
    and g1154 ( n11720 , n16767 , n4704 );
    not g1155 ( n1710 , n85 );
    or g1156 ( n28528 , n8100 , n22338 );
    or g1157 ( n25816 , n17305 , n21954 );
    or g1158 ( n2999 , n13640 , n25688 );
    xnor g1159 ( n6131 , n4277 , n7354 );
    xnor g1160 ( n7871 , n22104 , n31326 );
    and g1161 ( n23029 , n9828 , n16966 );
    not g1162 ( n460 , n15517 );
    or g1163 ( n13284 , n553 , n6370 );
    xnor g1164 ( n11612 , n5654 , n31970 );
    or g1165 ( n28184 , n15628 , n29701 );
    not g1166 ( n20779 , n28021 );
    and g1167 ( n18973 , n802 , n20517 );
    nor g1168 ( n1116 , n9146 , n21716 );
    not g1169 ( n23088 , n4934 );
    and g1170 ( n20047 , n11567 , n3003 );
    xnor g1171 ( n24725 , n2402 , n1964 );
    xor g1172 ( n29811 , n1091 , n18344 );
    not g1173 ( n27925 , n4728 );
    and g1174 ( n715 , n27436 , n1558 );
    nor g1175 ( n1764 , n2653 , n13485 );
    not g1176 ( n21114 , n4243 );
    not g1177 ( n14362 , n24086 );
    and g1178 ( n6662 , n4206 , n6998 );
    or g1179 ( n26528 , n25010 , n16897 );
    xor g1180 ( n27016 , n29202 , n10037 );
    not g1181 ( n10450 , n8873 );
    not g1182 ( n231 , n13405 );
    and g1183 ( n27697 , n23473 , n2837 );
    xnor g1184 ( n30969 , n20420 , n22746 );
    xnor g1185 ( n18817 , n11874 , n26029 );
    nor g1186 ( n12244 , n2629 , n17440 );
    or g1187 ( n8599 , n4798 , n21062 );
    nor g1188 ( n15796 , n17798 , n8572 );
    xnor g1189 ( n29388 , n15436 , n18551 );
    xnor g1190 ( n8384 , n29506 , n2675 );
    not g1191 ( n15109 , n16254 );
    nor g1192 ( n14680 , n21136 , n19217 );
    buf g1193 ( n23138 , n18035 );
    xnor g1194 ( n19295 , n19351 , n3287 );
    xor g1195 ( n5812 , n20533 , n23770 );
    nor g1196 ( n9044 , n26894 , n17843 );
    not g1197 ( n12112 , n24712 );
    not g1198 ( n10238 , n8865 );
    and g1199 ( n2117 , n5242 , n11841 );
    xnor g1200 ( n18856 , n13668 , n4358 );
    xnor g1201 ( n21216 , n890 , n4114 );
    or g1202 ( n24665 , n29732 , n17782 );
    not g1203 ( n6763 , n20134 );
    or g1204 ( n31036 , n13305 , n1142 );
    and g1205 ( n14927 , n23622 , n15291 );
    and g1206 ( n3161 , n30443 , n29700 );
    not g1207 ( n21676 , n18507 );
    not g1208 ( n3050 , n30817 );
    or g1209 ( n23211 , n8183 , n13265 );
    not g1210 ( n17579 , n8803 );
    and g1211 ( n7257 , n29585 , n11158 );
    or g1212 ( n13818 , n13350 , n31038 );
    nor g1213 ( n18565 , n6127 , n14499 );
    and g1214 ( n2843 , n23423 , n17759 );
    not g1215 ( n5708 , n29348 );
    or g1216 ( n26307 , n12803 , n10658 );
    not g1217 ( n8018 , n7336 );
    xnor g1218 ( n9388 , n866 , n6477 );
    xnor g1219 ( n19902 , n13862 , n20097 );
    xnor g1220 ( n25828 , n23482 , n1261 );
    xnor g1221 ( n12015 , n19409 , n10327 );
    and g1222 ( n4381 , n25634 , n6294 );
    nor g1223 ( n6870 , n10196 , n9029 );
    nor g1224 ( n30166 , n28973 , n5572 );
    not g1225 ( n26419 , n26131 );
    or g1226 ( n9692 , n15009 , n28968 );
    or g1227 ( n30976 , n1457 , n1298 );
    or g1228 ( n30007 , n5583 , n6175 );
    or g1229 ( n6045 , n23232 , n7086 );
    not g1230 ( n13191 , n21253 );
    or g1231 ( n8192 , n20291 , n30795 );
    or g1232 ( n25440 , n9483 , n5426 );
    or g1233 ( n11669 , n4065 , n2272 );
    not g1234 ( n27087 , n13754 );
    not g1235 ( n31806 , n22936 );
    not g1236 ( n12872 , n3475 );
    not g1237 ( n9189 , n15396 );
    not g1238 ( n15179 , n23444 );
    not g1239 ( n23693 , n554 );
    not g1240 ( n23099 , n15749 );
    buf g1241 ( n22746 , n15041 );
    nor g1242 ( n1538 , n8553 , n4160 );
    or g1243 ( n4055 , n8078 , n7328 );
    xnor g1244 ( n18823 , n20046 , n13543 );
    xnor g1245 ( n25391 , n6865 , n19222 );
    nor g1246 ( n25574 , n26117 , n3789 );
    xnor g1247 ( n9587 , n949 , n27403 );
    xnor g1248 ( n30347 , n5572 , n27948 );
    not g1249 ( n20691 , n22235 );
    xnor g1250 ( n22187 , n28507 , n28151 );
    or g1251 ( n2662 , n24371 , n17005 );
    or g1252 ( n13611 , n13566 , n31726 );
    not g1253 ( n18720 , n19600 );
    xnor g1254 ( n4034 , n15442 , n13826 );
    or g1255 ( n21623 , n14616 , n12156 );
    xnor g1256 ( n27792 , n4111 , n16891 );
    or g1257 ( n24042 , n15616 , n12787 );
    or g1258 ( n2905 , n29670 , n19963 );
    or g1259 ( n21121 , n1788 , n25941 );
    xnor g1260 ( n23248 , n30228 , n24929 );
    and g1261 ( n22320 , n26727 , n22862 );
    and g1262 ( n17546 , n2487 , n16056 );
    and g1263 ( n13349 , n27482 , n15258 );
    not g1264 ( n27218 , n13137 );
    not g1265 ( n8049 , n22688 );
    nor g1266 ( n14157 , n775 , n26148 );
    xnor g1267 ( n15079 , n21319 , n1539 );
    xnor g1268 ( n21220 , n10601 , n11223 );
    buf g1269 ( n30022 , n17195 );
    or g1270 ( n29760 , n29047 , n9878 );
    not g1271 ( n4500 , n28884 );
    xnor g1272 ( n6108 , n5904 , n24609 );
    xnor g1273 ( n24032 , n229 , n25807 );
    xnor g1274 ( n17919 , n1978 , n1345 );
    nor g1275 ( n14313 , n27638 , n22039 );
    xnor g1276 ( n24812 , n25727 , n11789 );
    xnor g1277 ( n29949 , n20317 , n7434 );
    xnor g1278 ( n26566 , n2328 , n9479 );
    not g1279 ( n14974 , n19512 );
    and g1280 ( n19579 , n25314 , n647 );
    xnor g1281 ( n14938 , n27526 , n31030 );
    xnor g1282 ( n19220 , n13882 , n11945 );
    or g1283 ( n5921 , n18355 , n27482 );
    or g1284 ( n22070 , n26879 , n9728 );
    xor g1285 ( n1717 , n30000 , n5948 );
    nor g1286 ( n16215 , n31111 , n3611 );
    not g1287 ( n23236 , n31191 );
    or g1288 ( n18273 , n31769 , n8557 );
    or g1289 ( n23908 , n4609 , n28690 );
    not g1290 ( n25958 , n14268 );
    not g1291 ( n30565 , n10139 );
    or g1292 ( n12006 , n1812 , n12034 );
    or g1293 ( n16447 , n6529 , n12040 );
    not g1294 ( n17812 , n21266 );
    not g1295 ( n25608 , n30775 );
    and g1296 ( n15958 , n21936 , n8564 );
    xnor g1297 ( n579 , n6744 , n14918 );
    or g1298 ( n3737 , n6243 , n25728 );
    not g1299 ( n5038 , n6883 );
    nor g1300 ( n9846 , n24429 , n13949 );
    or g1301 ( n28273 , n18243 , n13682 );
    and g1302 ( n9801 , n14120 , n2413 );
    not g1303 ( n12569 , n11561 );
    xnor g1304 ( n9724 , n17735 , n29452 );
    or g1305 ( n12085 , n9787 , n4502 );
    or g1306 ( n14933 , n17593 , n17549 );
    or g1307 ( n2114 , n25474 , n5278 );
    or g1308 ( n26405 , n25180 , n25088 );
    xnor g1309 ( n3576 , n30045 , n22922 );
    nor g1310 ( n5376 , n27196 , n15470 );
    not g1311 ( n29581 , n30649 );
    nor g1312 ( n9265 , n11232 , n19432 );
    not g1313 ( n15429 , n9885 );
    xnor g1314 ( n8632 , n21050 , n26894 );
    and g1315 ( n4636 , n12227 , n5127 );
    not g1316 ( n2019 , n18707 );
    xnor g1317 ( n20214 , n18246 , n11601 );
    not g1318 ( n4248 , n7122 );
    and g1319 ( n10437 , n4024 , n31991 );
    not g1320 ( n8862 , n4868 );
    and g1321 ( n25593 , n2387 , n11336 );
    xnor g1322 ( n1242 , n1616 , n3036 );
    xnor g1323 ( n19706 , n30635 , n803 );
    xnor g1324 ( n31955 , n8409 , n9058 );
    xnor g1325 ( n15494 , n7326 , n16714 );
    not g1326 ( n7090 , n31979 );
    xnor g1327 ( n23703 , n31931 , n983 );
    not g1328 ( n30746 , n29978 );
    and g1329 ( n31861 , n9085 , n2142 );
    not g1330 ( n8361 , n1935 );
    not g1331 ( n27074 , n18096 );
    not g1332 ( n9373 , n9071 );
    or g1333 ( n24470 , n1505 , n24778 );
    nor g1334 ( n6648 , n8986 , n31889 );
    not g1335 ( n5274 , n5030 );
    xnor g1336 ( n17872 , n9655 , n24429 );
    or g1337 ( n3504 , n13738 , n15282 );
    xnor g1338 ( n29310 , n2690 , n22675 );
    xnor g1339 ( n30692 , n19922 , n29520 );
    or g1340 ( n26621 , n5930 , n4433 );
    or g1341 ( n21247 , n6568 , n23809 );
    not g1342 ( n5342 , n22866 );
    or g1343 ( n2279 , n7091 , n21898 );
    xnor g1344 ( n4642 , n31680 , n26836 );
    xor g1345 ( n21063 , n23632 , n664 );
    not g1346 ( n15711 , n13405 );
    not g1347 ( n7229 , n11736 );
    or g1348 ( n9704 , n28648 , n11690 );
    nor g1349 ( n27612 , n8312 , n16882 );
    not g1350 ( n2238 , n9970 );
    and g1351 ( n15885 , n23500 , n1009 );
    xnor g1352 ( n5544 , n27126 , n9424 );
    and g1353 ( n13902 , n15929 , n21708 );
    or g1354 ( n30134 , n3502 , n28883 );
    xnor g1355 ( n19878 , n21032 , n19394 );
    and g1356 ( n21550 , n13231 , n21254 );
    xnor g1357 ( n13018 , n16411 , n12566 );
    not g1358 ( n24195 , n26799 );
    or g1359 ( n22653 , n14633 , n22795 );
    buf g1360 ( n12221 , n21684 );
    not g1361 ( n24704 , n21485 );
    xnor g1362 ( n4720 , n17417 , n26961 );
    or g1363 ( n17577 , n18388 , n19101 );
    not g1364 ( n23223 , n9469 );
    xnor g1365 ( n8780 , n15023 , n3418 );
    xnor g1366 ( n26512 , n26281 , n7315 );
    xnor g1367 ( n22530 , n7515 , n29947 );
    or g1368 ( n44 , n25192 , n21072 );
    not g1369 ( n1192 , n30453 );
    xnor g1370 ( n26606 , n7172 , n7900 );
    xnor g1371 ( n23411 , n20495 , n16609 );
    xnor g1372 ( n27502 , n13881 , n21672 );
    not g1373 ( n12396 , n29390 );
    xnor g1374 ( n1727 , n21172 , n23996 );
    xnor g1375 ( n25331 , n4229 , n6230 );
    or g1376 ( n15302 , n21276 , n2256 );
    or g1377 ( n31347 , n10499 , n16802 );
    and g1378 ( n16446 , n8605 , n7780 );
    not g1379 ( n27597 , n1427 );
    xnor g1380 ( n5256 , n13363 , n1354 );
    not g1381 ( n26675 , n18118 );
    not g1382 ( n27175 , n25857 );
    nor g1383 ( n17556 , n7933 , n4370 );
    not g1384 ( n24735 , n29857 );
    xnor g1385 ( n2240 , n3311 , n124 );
    or g1386 ( n2101 , n6016 , n10997 );
    nor g1387 ( n15699 , n14956 , n10040 );
    xnor g1388 ( n30386 , n16160 , n14470 );
    xnor g1389 ( n1301 , n22976 , n28654 );
    or g1390 ( n22278 , n1616 , n10302 );
    and g1391 ( n130 , n3697 , n17017 );
    xnor g1392 ( n3526 , n25118 , n28432 );
    xnor g1393 ( n13404 , n23184 , n1518 );
    or g1394 ( n5818 , n3690 , n23704 );
    and g1395 ( n21976 , n6899 , n7519 );
    or g1396 ( n16726 , n13680 , n17833 );
    or g1397 ( n24119 , n19025 , n21561 );
    or g1398 ( n21440 , n17733 , n6851 );
    not g1399 ( n2383 , n7141 );
    or g1400 ( n10188 , n11805 , n17458 );
    not g1401 ( n5786 , n4831 );
    or g1402 ( n30032 , n9019 , n12644 );
    or g1403 ( n19470 , n19757 , n13896 );
    nor g1404 ( n12326 , n14680 , n22630 );
    xnor g1405 ( n24487 , n22051 , n9228 );
    not g1406 ( n1058 , n27578 );
    xnor g1407 ( n17776 , n2169 , n13834 );
    not g1408 ( n22028 , n3996 );
    or g1409 ( n29565 , n29958 , n18944 );
    and g1410 ( n21924 , n31887 , n218 );
    and g1411 ( n9932 , n31678 , n2333 );
    not g1412 ( n546 , n7021 );
    and g1413 ( n25343 , n17137 , n25552 );
    and g1414 ( n7018 , n27249 , n21433 );
    nor g1415 ( n11599 , n1705 , n31958 );
    xnor g1416 ( n22236 , n7213 , n22607 );
    and g1417 ( n6452 , n7421 , n7900 );
    not g1418 ( n22815 , n4624 );
    xnor g1419 ( n8771 , n29735 , n14668 );
    xnor g1420 ( n24848 , n22867 , n24429 );
    xnor g1421 ( n11963 , n15032 , n13961 );
    xnor g1422 ( n27937 , n28951 , n2629 );
    nor g1423 ( n28193 , n14992 , n21824 );
    xnor g1424 ( n17163 , n14227 , n13526 );
    nor g1425 ( n2912 , n25305 , n21720 );
    or g1426 ( n4357 , n15213 , n22004 );
    not g1427 ( n27430 , n21841 );
    nor g1428 ( n1850 , n9469 , n25904 );
    nor g1429 ( n18819 , n10474 , n31847 );
    or g1430 ( n31771 , n2787 , n3805 );
    nor g1431 ( n15135 , n23172 , n3784 );
    not g1432 ( n798 , n17255 );
    or g1433 ( n23007 , n25635 , n6884 );
    nor g1434 ( n21140 , n13764 , n8915 );
    xnor g1435 ( n23844 , n3497 , n25498 );
    xnor g1436 ( n15951 , n3941 , n9837 );
    or g1437 ( n22416 , n5126 , n833 );
    nor g1438 ( n8006 , n24129 , n26346 );
    not g1439 ( n16340 , n445 );
    xnor g1440 ( n10408 , n11024 , n1481 );
    not g1441 ( n24386 , n11642 );
    not g1442 ( n18604 , n7216 );
    or g1443 ( n8684 , n3382 , n16175 );
    not g1444 ( n20525 , n31965 );
    or g1445 ( n703 , n25577 , n19400 );
    and g1446 ( n10116 , n25468 , n19772 );
    not g1447 ( n24875 , n13943 );
    not g1448 ( n5609 , n10730 );
    and g1449 ( n19553 , n19154 , n8840 );
    not g1450 ( n16740 , n8622 );
    and g1451 ( n9192 , n28799 , n28749 );
    not g1452 ( n9996 , n19189 );
    nor g1453 ( n23446 , n23557 , n29163 );
    and g1454 ( n29850 , n26586 , n3510 );
    or g1455 ( n15647 , n12181 , n31288 );
    xnor g1456 ( n21204 , n1480 , n13094 );
    or g1457 ( n7961 , n9800 , n28492 );
    or g1458 ( n12422 , n14719 , n23543 );
    not g1459 ( n10243 , n27555 );
    and g1460 ( n31439 , n8813 , n21994 );
    not g1461 ( n20086 , n18551 );
    or g1462 ( n12973 , n11189 , n15685 );
    xnor g1463 ( n10019 , n23452 , n21895 );
    not g1464 ( n19036 , n17801 );
    or g1465 ( n32030 , n17136 , n25831 );
    nor g1466 ( n24730 , n4696 , n8357 );
    or g1467 ( n31531 , n9711 , n20071 );
    xnor g1468 ( n23552 , n19102 , n12607 );
    and g1469 ( n22689 , n28466 , n10237 );
    xnor g1470 ( n4214 , n10432 , n30831 );
    not g1471 ( n215 , n9933 );
    and g1472 ( n31422 , n15450 , n12403 );
    and g1473 ( n22067 , n7985 , n11403 );
    xnor g1474 ( n31863 , n19357 , n25798 );
    xnor g1475 ( n20304 , n4186 , n25476 );
    xor g1476 ( n26940 , n2609 , n28801 );
    or g1477 ( n27136 , n4668 , n11960 );
    or g1478 ( n10436 , n28594 , n4378 );
    xnor g1479 ( n20504 , n29178 , n16278 );
    or g1480 ( n12163 , n4192 , n25136 );
    xnor g1481 ( n14063 , n1583 , n17119 );
    or g1482 ( n25270 , n24234 , n3247 );
    or g1483 ( n28344 , n25024 , n22072 );
    not g1484 ( n4074 , n5174 );
    not g1485 ( n2792 , n29617 );
    nor g1486 ( n29283 , n20482 , n5500 );
    and g1487 ( n3277 , n9843 , n1819 );
    xnor g1488 ( n29744 , n25527 , n27453 );
    not g1489 ( n30024 , n20788 );
    not g1490 ( n28683 , n170 );
    not g1491 ( n5984 , n4075 );
    nor g1492 ( n21078 , n4264 , n24236 );
    not g1493 ( n29414 , n22886 );
    and g1494 ( n28744 , n5849 , n7153 );
    not g1495 ( n11644 , n8960 );
    not g1496 ( n7055 , n18380 );
    not g1497 ( n29066 , n13196 );
    nor g1498 ( n12763 , n21009 , n27570 );
    not g1499 ( n14422 , n20100 );
    not g1500 ( n8929 , n10689 );
    and g1501 ( n31825 , n10164 , n14254 );
    or g1502 ( n17647 , n27891 , n6232 );
    xnor g1503 ( n11353 , n8224 , n25048 );
    not g1504 ( n29978 , n11323 );
    xnor g1505 ( n18244 , n18483 , n288 );
    and g1506 ( n14414 , n11533 , n30669 );
    nor g1507 ( n20833 , n6127 , n6787 );
    or g1508 ( n1834 , n2877 , n25051 );
    not g1509 ( n31989 , n14380 );
    xnor g1510 ( n19388 , n27075 , n15987 );
    nor g1511 ( n19450 , n14424 , n17893 );
    xnor g1512 ( n6330 , n30365 , n8046 );
    or g1513 ( n27333 , n10433 , n10598 );
    xnor g1514 ( n3752 , n22630 , n27754 );
    or g1515 ( n18634 , n18925 , n27389 );
    not g1516 ( n3408 , n2864 );
    xnor g1517 ( n10088 , n7116 , n892 );
    nor g1518 ( n28757 , n15178 , n7701 );
    or g1519 ( n28846 , n15259 , n9700 );
    not g1520 ( n1188 , n22803 );
    and g1521 ( n6020 , n7149 , n16532 );
    and g1522 ( n29999 , n27591 , n22423 );
    not g1523 ( n10479 , n5569 );
    nor g1524 ( n10721 , n21133 , n1072 );
    nor g1525 ( n10421 , n19134 , n316 );
    nor g1526 ( n17013 , n2283 , n28068 );
    xor g1527 ( n2491 , n18873 , n1653 );
    xnor g1528 ( n19796 , n26099 , n27274 );
    not g1529 ( n11082 , n4790 );
    xnor g1530 ( n22827 , n30418 , n6874 );
    not g1531 ( n30945 , n10015 );
    or g1532 ( n15046 , n15912 , n28148 );
    or g1533 ( n19627 , n16917 , n7716 );
    xnor g1534 ( n29559 , n21704 , n29682 );
    or g1535 ( n4203 , n8808 , n3600 );
    and g1536 ( n2622 , n29555 , n9153 );
    not g1537 ( n1570 , n21928 );
    xnor g1538 ( n15148 , n8651 , n9545 );
    nor g1539 ( n3554 , n19597 , n11856 );
    or g1540 ( n18130 , n5336 , n31271 );
    xnor g1541 ( n9888 , n9042 , n1126 );
    xnor g1542 ( n6174 , n18497 , n488 );
    xnor g1543 ( n15115 , n3020 , n16146 );
    and g1544 ( n15923 , n30714 , n27856 );
    and g1545 ( n9698 , n3421 , n13777 );
    or g1546 ( n7383 , n23715 , n14378 );
    not g1547 ( n17514 , n14946 );
    or g1548 ( n15057 , n18712 , n26169 );
    and g1549 ( n25943 , n13136 , n22927 );
    nor g1550 ( n549 , n21064 , n26866 );
    and g1551 ( n3798 , n3589 , n27594 );
    not g1552 ( n12186 , n30793 );
    or g1553 ( n6102 , n24455 , n19101 );
    not g1554 ( n12067 , n8451 );
    or g1555 ( n11661 , n2176 , n30482 );
    not g1556 ( n2628 , n4213 );
    not g1557 ( n10895 , n27354 );
    or g1558 ( n17175 , n8360 , n31976 );
    nor g1559 ( n24757 , n20067 , n24935 );
    or g1560 ( n23055 , n27948 , n27129 );
    not g1561 ( n30369 , n13869 );
    and g1562 ( n6397 , n11181 , n16168 );
    and g1563 ( n13927 , n19409 , n25851 );
    not g1564 ( n29895 , n19420 );
    and g1565 ( n29651 , n15984 , n8892 );
    xnor g1566 ( n22620 , n11559 , n8754 );
    or g1567 ( n9686 , n26306 , n21964 );
    or g1568 ( n9510 , n12932 , n13207 );
    xnor g1569 ( n8240 , n17030 , n8988 );
    xnor g1570 ( n10204 , n23207 , n11215 );
    not g1571 ( n10926 , n17844 );
    nor g1572 ( n5434 , n19615 , n14999 );
    or g1573 ( n25770 , n23008 , n733 );
    and g1574 ( n28886 , n3061 , n15486 );
    not g1575 ( n29839 , n14965 );
    or g1576 ( n1298 , n709 , n28275 );
    and g1577 ( n27066 , n2131 , n15066 );
    or g1578 ( n4808 , n26191 , n22528 );
    nor g1579 ( n11195 , n22045 , n18380 );
    or g1580 ( n1395 , n21789 , n20652 );
    nor g1581 ( n14094 , n9626 , n25012 );
    or g1582 ( n19827 , n13718 , n11359 );
    xnor g1583 ( n31440 , n2154 , n6927 );
    and g1584 ( n25401 , n7628 , n20540 );
    or g1585 ( n29489 , n24661 , n12894 );
    nor g1586 ( n12874 , n5149 , n12771 );
    nor g1587 ( n12989 , n29695 , n16723 );
    xnor g1588 ( n23828 , n20893 , n17147 );
    and g1589 ( n1311 , n22065 , n16773 );
    and g1590 ( n12563 , n31361 , n13725 );
    or g1591 ( n31065 , n7493 , n15116 );
    not g1592 ( n16255 , n26469 );
    or g1593 ( n24799 , n27149 , n28002 );
    not g1594 ( n9925 , n2978 );
    xnor g1595 ( n31281 , n1947 , n169 );
    xnor g1596 ( n11307 , n14651 , n2732 );
    xnor g1597 ( n26266 , n9589 , n30457 );
    not g1598 ( n20897 , n15991 );
    not g1599 ( n13506 , n4484 );
    and g1600 ( n27858 , n2366 , n5445 );
    xnor g1601 ( n5095 , n10391 , n4165 );
    xnor g1602 ( n870 , n23063 , n15126 );
    xnor g1603 ( n17367 , n908 , n8987 );
    not g1604 ( n25042 , n18227 );
    not g1605 ( n22610 , n5901 );
    xnor g1606 ( n11498 , n19480 , n14917 );
    xnor g1607 ( n14231 , n24423 , n2438 );
    or g1608 ( n18220 , n28645 , n19672 );
    not g1609 ( n4592 , n6052 );
    xnor g1610 ( n23666 , n29799 , n4368 );
    and g1611 ( n20321 , n2257 , n26291 );
    or g1612 ( n4139 , n21786 , n20476 );
    xor g1613 ( n7323 , n19786 , n30826 );
    or g1614 ( n12107 , n31471 , n6875 );
    or g1615 ( n5705 , n5784 , n29438 );
    or g1616 ( n16346 , n818 , n9026 );
    and g1617 ( n741 , n5894 , n23804 );
    or g1618 ( n691 , n5607 , n19669 );
    xnor g1619 ( n31831 , n6113 , n15300 );
    and g1620 ( n29515 , n21304 , n22376 );
    or g1621 ( n20619 , n21180 , n5159 );
    and g1622 ( n1016 , n26668 , n13707 );
    and g1623 ( n17229 , n26265 , n3432 );
    or g1624 ( n18046 , n14168 , n17690 );
    xnor g1625 ( n14913 , n2875 , n9904 );
    nor g1626 ( n25158 , n4674 , n4294 );
    or g1627 ( n27480 , n6053 , n5613 );
    not g1628 ( n32010 , n31800 );
    or g1629 ( n29864 , n7035 , n30015 );
    xnor g1630 ( n31210 , n15663 , n3591 );
    xnor g1631 ( n14870 , n7636 , n21381 );
    or g1632 ( n21189 , n8985 , n2773 );
    nor g1633 ( n13226 , n13194 , n12425 );
    and g1634 ( n23080 , n1209 , n27485 );
    or g1635 ( n3533 , n31896 , n14104 );
    xnor g1636 ( n26817 , n18302 , n15283 );
    nor g1637 ( n19495 , n25649 , n12226 );
    not g1638 ( n12333 , n25987 );
    nor g1639 ( n12515 , n643 , n10882 );
    and g1640 ( n2376 , n7888 , n23376 );
    or g1641 ( n913 , n1953 , n4065 );
    xnor g1642 ( n19261 , n2363 , n5915 );
    nor g1643 ( n8131 , n32002 , n9989 );
    and g1644 ( n25418 , n1070 , n12855 );
    or g1645 ( n6899 , n21960 , n31586 );
    xnor g1646 ( n12707 , n14551 , n3285 );
    xnor g1647 ( n9302 , n17318 , n29368 );
    not g1648 ( n742 , n5172 );
    and g1649 ( n9826 , n30995 , n8280 );
    xnor g1650 ( n1529 , n19950 , n27940 );
    not g1651 ( n15939 , n29129 );
    or g1652 ( n4853 , n25062 , n849 );
    not g1653 ( n14843 , n30808 );
    or g1654 ( n29154 , n29151 , n26738 );
    not g1655 ( n13682 , n15105 );
    not g1656 ( n21984 , n19059 );
    not g1657 ( n12367 , n18165 );
    xnor g1658 ( n24743 , n28417 , n350 );
    xnor g1659 ( n29105 , n12820 , n5546 );
    and g1660 ( n22101 , n27468 , n15250 );
    not g1661 ( n31391 , n14366 );
    not g1662 ( n18520 , n6756 );
    xor g1663 ( n7381 , n9814 , n17505 );
    xnor g1664 ( n31197 , n19208 , n16117 );
    xnor g1665 ( n7788 , n19373 , n21485 );
    not g1666 ( n9832 , n3283 );
    or g1667 ( n18638 , n17267 , n3008 );
    and g1668 ( n26275 , n704 , n25334 );
    not g1669 ( n26605 , n1040 );
    and g1670 ( n1631 , n24460 , n11165 );
    and g1671 ( n10984 , n24922 , n10694 );
    nor g1672 ( n26369 , n22366 , n4227 );
    not g1673 ( n3401 , n18139 );
    not g1674 ( n17664 , n19861 );
    xnor g1675 ( n28945 , n7449 , n12751 );
    not g1676 ( n12883 , n18751 );
    nor g1677 ( n6093 , n7655 , n27430 );
    nor g1678 ( n24334 , n14356 , n2395 );
    or g1679 ( n4971 , n21896 , n1557 );
    not g1680 ( n2222 , n10742 );
    not g1681 ( n26568 , n23963 );
    or g1682 ( n18001 , n17227 , n27885 );
    xnor g1683 ( n27657 , n22708 , n30529 );
    not g1684 ( n12837 , n5300 );
    xnor g1685 ( n6338 , n18123 , n25920 );
    or g1686 ( n20972 , n27653 , n15062 );
    xnor g1687 ( n25133 , n24468 , n8183 );
    and g1688 ( n1975 , n18911 , n3583 );
    xnor g1689 ( n25329 , n4998 , n18608 );
    or g1690 ( n16336 , n27606 , n4660 );
    and g1691 ( n24854 , n3901 , n13806 );
    xnor g1692 ( n8515 , n23810 , n3034 );
    or g1693 ( n6869 , n27586 , n5421 );
    or g1694 ( n28415 , n18148 , n25164 );
    not g1695 ( n240 , n23907 );
    xnor g1696 ( n1042 , n29019 , n26002 );
    xnor g1697 ( n24107 , n22922 , n24066 );
    not g1698 ( n24136 , n28045 );
    not g1699 ( n22570 , n12488 );
    xnor g1700 ( n5341 , n12917 , n30 );
    and g1701 ( n2601 , n3151 , n29941 );
    xnor g1702 ( n21722 , n16823 , n10680 );
    xnor g1703 ( n15174 , n179 , n344 );
    or g1704 ( n29221 , n26514 , n382 );
    nor g1705 ( n14072 , n20198 , n23437 );
    or g1706 ( n12752 , n5134 , n16073 );
    not g1707 ( n2975 , n7710 );
    not g1708 ( n21058 , n23828 );
    or g1709 ( n26638 , n26440 , n25743 );
    and g1710 ( n6678 , n2045 , n14071 );
    or g1711 ( n6190 , n4205 , n17956 );
    xnor g1712 ( n7267 , n13639 , n27442 );
    not g1713 ( n15721 , n18897 );
    or g1714 ( n5186 , n26897 , n30946 );
    nor g1715 ( n27586 , n10393 , n27121 );
    xnor g1716 ( n15927 , n10416 , n6560 );
    not g1717 ( n1900 , n4512 );
    or g1718 ( n27909 , n23941 , n7770 );
    nor g1719 ( n25084 , n10363 , n14711 );
    not g1720 ( n18344 , n2337 );
    not g1721 ( n14597 , n6541 );
    not g1722 ( n23761 , n19254 );
    not g1723 ( n17652 , n5272 );
    xnor g1724 ( n11233 , n11927 , n24940 );
    not g1725 ( n11211 , n7561 );
    or g1726 ( n28560 , n25099 , n22669 );
    not g1727 ( n13600 , n28614 );
    not g1728 ( n2259 , n5880 );
    or g1729 ( n26441 , n5984 , n11110 );
    xnor g1730 ( n29196 , n9950 , n8324 );
    or g1731 ( n12850 , n19940 , n12361 );
    xnor g1732 ( n2346 , n5433 , n3877 );
    not g1733 ( n1487 , n6937 );
    not g1734 ( n1705 , n8844 );
    or g1735 ( n10298 , n24532 , n4671 );
    or g1736 ( n11219 , n14242 , n25573 );
    not g1737 ( n27731 , n7705 );
    and g1738 ( n27170 , n17231 , n22523 );
    nor g1739 ( n20666 , n2248 , n257 );
    xnor g1740 ( n17375 , n22422 , n23047 );
    or g1741 ( n4741 , n15957 , n1544 );
    xnor g1742 ( n10724 , n9757 , n1767 );
    nor g1743 ( n9544 , n18391 , n9619 );
    nor g1744 ( n22963 , n16785 , n22934 );
    xnor g1745 ( n6105 , n20207 , n30064 );
    xnor g1746 ( n10475 , n11882 , n8466 );
    nor g1747 ( n5755 , n2444 , n22870 );
    and g1748 ( n31906 , n19832 , n15568 );
    or g1749 ( n19606 , n5540 , n24009 );
    xnor g1750 ( n27750 , n1348 , n17927 );
    nor g1751 ( n10331 , n7147 , n22708 );
    nor g1752 ( n5492 , n19231 , n12694 );
    or g1753 ( n25582 , n25897 , n14042 );
    or g1754 ( n14759 , n30291 , n4416 );
    and g1755 ( n20863 , n29658 , n12929 );
    not g1756 ( n12730 , n27235 );
    and g1757 ( n9571 , n5975 , n4168 );
    or g1758 ( n5748 , n15713 , n20985 );
    not g1759 ( n30102 , n1997 );
    xnor g1760 ( n30009 , n17185 , n6895 );
    xnor g1761 ( n4027 , n18389 , n13526 );
    or g1762 ( n22171 , n14406 , n24764 );
    xnor g1763 ( n21188 , n25055 , n18846 );
    not g1764 ( n7131 , n24363 );
    or g1765 ( n10079 , n23185 , n2990 );
    not g1766 ( n12618 , n23490 );
    xnor g1767 ( n21073 , n10433 , n23115 );
    and g1768 ( n6575 , n3598 , n28457 );
    or g1769 ( n26411 , n9370 , n5898 );
    not g1770 ( n29134 , n508 );
    not g1771 ( n29199 , n28210 );
    xnor g1772 ( n8820 , n9899 , n6963 );
    and g1773 ( n13396 , n10103 , n16808 );
    and g1774 ( n21388 , n14877 , n22784 );
    buf g1775 ( n2753 , n29963 );
    and g1776 ( n12101 , n26581 , n12935 );
    xnor g1777 ( n30930 , n22273 , n12462 );
    and g1778 ( n24084 , n14648 , n14992 );
    or g1779 ( n18405 , n595 , n14426 );
    xnor g1780 ( n26880 , n25944 , n26914 );
    or g1781 ( n17091 , n4667 , n5286 );
    and g1782 ( n13282 , n1938 , n472 );
    not g1783 ( n8241 , n26306 );
    and g1784 ( n23216 , n22011 , n7030 );
    xor g1785 ( n7216 , n25548 , n14690 );
    not g1786 ( n19728 , n3021 );
    xnor g1787 ( n10375 , n16772 , n21493 );
    or g1788 ( n23442 , n27242 , n19428 );
    xnor g1789 ( n8125 , n26304 , n31624 );
    not g1790 ( n8300 , n16676 );
    xnor g1791 ( n26751 , n31253 , n8168 );
    not g1792 ( n13032 , n14328 );
    or g1793 ( n27548 , n24485 , n8661 );
    nor g1794 ( n27079 , n18095 , n10683 );
    not g1795 ( n5991 , n16128 );
    or g1796 ( n17671 , n3771 , n1336 );
    and g1797 ( n25139 , n17770 , n11664 );
    not g1798 ( n13279 , n13271 );
    nor g1799 ( n27462 , n23163 , n21198 );
    not g1800 ( n220 , n19593 );
    or g1801 ( n8353 , n3591 , n31091 );
    or g1802 ( n20581 , n27799 , n26874 );
    xnor g1803 ( n4529 , n6059 , n22007 );
    and g1804 ( n6091 , n24686 , n14497 );
    xnor g1805 ( n7747 , n21450 , n13939 );
    xnor g1806 ( n23461 , n750 , n3511 );
    or g1807 ( n10672 , n29723 , n8420 );
    xnor g1808 ( n2949 , n18376 , n29604 );
    or g1809 ( n19195 , n25567 , n3684 );
    nor g1810 ( n867 , n24132 , n23400 );
    xnor g1811 ( n14081 , n29075 , n30505 );
    xnor g1812 ( n27940 , n10047 , n1995 );
    and g1813 ( n15675 , n23030 , n22290 );
    or g1814 ( n19964 , n4175 , n26695 );
    or g1815 ( n27240 , n22560 , n6370 );
    or g1816 ( n16971 , n12028 , n12971 );
    and g1817 ( n17569 , n24267 , n29379 );
    not g1818 ( n11800 , n30873 );
    and g1819 ( n2967 , n26722 , n6028 );
    and g1820 ( n268 , n6582 , n21788 );
    xnor g1821 ( n29474 , n4024 , n16415 );
    not g1822 ( n20704 , n29084 );
    xnor g1823 ( n11209 , n22522 , n12207 );
    or g1824 ( n15051 , n3163 , n30370 );
    or g1825 ( n3790 , n21411 , n9913 );
    xnor g1826 ( n10653 , n5286 , n9659 );
    and g1827 ( n29919 , n23007 , n10632 );
    xnor g1828 ( n15487 , n14022 , n10961 );
    and g1829 ( n157 , n4117 , n20967 );
    not g1830 ( n2120 , n26354 );
    not g1831 ( n18243 , n17368 );
    xnor g1832 ( n15535 , n13872 , n2995 );
    or g1833 ( n29146 , n6773 , n24060 );
    xnor g1834 ( n21672 , n30429 , n11434 );
    and g1835 ( n16977 , n30563 , n29669 );
    or g1836 ( n24082 , n16344 , n28581 );
    not g1837 ( n12217 , n8563 );
    nor g1838 ( n25437 , n29185 , n19560 );
    not g1839 ( n26639 , n24429 );
    nor g1840 ( n16044 , n16474 , n1019 );
    xor g1841 ( n19158 , n9882 , n340 );
    not g1842 ( n2591 , n14894 );
    xnor g1843 ( n2404 , n5011 , n5265 );
    not g1844 ( n2814 , n22351 );
    not g1845 ( n27148 , n14421 );
    nor g1846 ( n25829 , n31316 , n30861 );
    xnor g1847 ( n15207 , n23481 , n17189 );
    not g1848 ( n1962 , n28856 );
    and g1849 ( n2664 , n29311 , n8751 );
    and g1850 ( n8024 , n14902 , n14196 );
    or g1851 ( n25631 , n14256 , n1438 );
    or g1852 ( n8066 , n8952 , n31997 );
    or g1853 ( n12391 , n6603 , n28857 );
    or g1854 ( n17685 , n31758 , n8866 );
    not g1855 ( n10466 , n12117 );
    not g1856 ( n7421 , n2127 );
    xnor g1857 ( n7075 , n3503 , n14479 );
    or g1858 ( n19795 , n5682 , n25250 );
    not g1859 ( n2428 , n21124 );
    and g1860 ( n29875 , n12249 , n216 );
    xnor g1861 ( n25267 , n1692 , n11643 );
    not g1862 ( n2026 , n17417 );
    and g1863 ( n14321 , n22684 , n20707 );
    nor g1864 ( n31241 , n31773 , n13510 );
    and g1865 ( n21571 , n23428 , n9891 );
    or g1866 ( n32031 , n25202 , n12091 );
    not g1867 ( n14940 , n7044 );
    xnor g1868 ( n22846 , n30313 , n30578 );
    not g1869 ( n5142 , n13970 );
    xnor g1870 ( n12717 , n21052 , n7589 );
    not g1871 ( n29681 , n18873 );
    or g1872 ( n3897 , n19779 , n24919 );
    or g1873 ( n23424 , n20132 , n16160 );
    and g1874 ( n23048 , n14840 , n9839 );
    not g1875 ( n18631 , n1453 );
    xor g1876 ( n23256 , n10960 , n9653 );
    or g1877 ( n16591 , n8970 , n29326 );
    xnor g1878 ( n3338 , n14169 , n14320 );
    not g1879 ( n10599 , n29982 );
    and g1880 ( n4790 , n11803 , n719 );
    or g1881 ( n7177 , n29355 , n1999 );
    not g1882 ( n1236 , n10355 );
    nor g1883 ( n612 , n10760 , n27490 );
    or g1884 ( n5658 , n26821 , n22975 );
    xnor g1885 ( n795 , n6881 , n7291 );
    or g1886 ( n22127 , n25127 , n11808 );
    not g1887 ( n9025 , n21447 );
    not g1888 ( n21928 , n4872 );
    not g1889 ( n26144 , n17079 );
    not g1890 ( n11104 , n28637 );
    not g1891 ( n17300 , n574 );
    and g1892 ( n27897 , n2831 , n9340 );
    not g1893 ( n5867 , n8475 );
    not g1894 ( n21988 , n5881 );
    or g1895 ( n29687 , n30342 , n21683 );
    not g1896 ( n30518 , n3884 );
    not g1897 ( n19529 , n29409 );
    xnor g1898 ( n1554 , n30238 , n20038 );
    not g1899 ( n19143 , n30085 );
    and g1900 ( n30807 , n9577 , n9522 );
    xnor g1901 ( n15914 , n28793 , n3392 );
    and g1902 ( n20512 , n1816 , n11282 );
    not g1903 ( n9830 , n10386 );
    not g1904 ( n4219 , n12079 );
    xnor g1905 ( n2034 , n29327 , n1700 );
    xnor g1906 ( n6453 , n8880 , n21949 );
    or g1907 ( n30267 , n19533 , n27346 );
    xnor g1908 ( n29021 , n13554 , n1980 );
    nor g1909 ( n26800 , n25452 , n28755 );
    or g1910 ( n6205 , n1039 , n4836 );
    not g1911 ( n14122 , n12035 );
    buf g1912 ( n20168 , n4326 );
    xnor g1913 ( n11071 , n20175 , n2825 );
    or g1914 ( n32026 , n7639 , n14568 );
    not g1915 ( n5494 , n27058 );
    xnor g1916 ( n30115 , n26736 , n12595 );
    not g1917 ( n24611 , n19937 );
    xnor g1918 ( n20665 , n8027 , n30031 );
    xnor g1919 ( n12096 , n29814 , n8393 );
    xnor g1920 ( n17830 , n13647 , n23476 );
    or g1921 ( n23500 , n5072 , n22239 );
    nor g1922 ( n4820 , n25265 , n11646 );
    and g1923 ( n7445 , n20577 , n12410 );
    nor g1924 ( n28700 , n27534 , n11537 );
    not g1925 ( n9575 , n27574 );
    not g1926 ( n1652 , n17151 );
    xnor g1927 ( n16561 , n18180 , n23346 );
    or g1928 ( n9160 , n18518 , n22659 );
    and g1929 ( n13487 , n2244 , n30961 );
    not g1930 ( n16930 , n6924 );
    xnor g1931 ( n3943 , n15003 , n14177 );
    not g1932 ( n4670 , n16558 );
    xnor g1933 ( n6686 , n5615 , n9075 );
    or g1934 ( n25878 , n3462 , n22650 );
    not g1935 ( n30180 , n21669 );
    and g1936 ( n28412 , n23872 , n20243 );
    or g1937 ( n30358 , n6193 , n30683 );
    and g1938 ( n16717 , n3219 , n28415 );
    not g1939 ( n2794 , n24429 );
    or g1940 ( n6155 , n1749 , n26059 );
    and g1941 ( n9770 , n27702 , n28086 );
    xnor g1942 ( n21468 , n22923 , n15220 );
    xnor g1943 ( n6369 , n19217 , n9653 );
    buf g1944 ( n13393 , n15891 );
    not g1945 ( n27216 , n7341 );
    and g1946 ( n31407 , n24762 , n25 );
    xnor g1947 ( n19251 , n9600 , n12663 );
    and g1948 ( n27490 , n17942 , n10121 );
    or g1949 ( n10885 , n2521 , n6560 );
    or g1950 ( n2707 , n29124 , n9771 );
    and g1951 ( n22765 , n29430 , n20536 );
    nor g1952 ( n2904 , n10139 , n31060 );
    not g1953 ( n19647 , n29647 );
    or g1954 ( n16635 , n23826 , n300 );
    not g1955 ( n14424 , n21246 );
    not g1956 ( n16105 , n16909 );
    not g1957 ( n14495 , n9163 );
    not g1958 ( n11641 , n20632 );
    or g1959 ( n20818 , n30152 , n14415 );
    not g1960 ( n15539 , n2791 );
    and g1961 ( n30883 , n31372 , n13552 );
    xnor g1962 ( n7632 , n893 , n8713 );
    not g1963 ( n25169 , n23158 );
    xnor g1964 ( n7755 , n4684 , n10014 );
    xnor g1965 ( n6054 , n28104 , n3113 );
    not g1966 ( n12410 , n27384 );
    or g1967 ( n25096 , n10433 , n18260 );
    nor g1968 ( n30193 , n10433 , n20289 );
    or g1969 ( n28354 , n31074 , n4995 );
    xnor g1970 ( n24513 , n9789 , n32007 );
    xnor g1971 ( n10569 , n14647 , n19162 );
    xnor g1972 ( n27898 , n25800 , n23653 );
    and g1973 ( n13446 , n2249 , n5094 );
    or g1974 ( n20932 , n28984 , n14853 );
    or g1975 ( n30524 , n13310 , n17654 );
    not g1976 ( n18355 , n13802 );
    xnor g1977 ( n28277 , n16076 , n7593 );
    xnor g1978 ( n7227 , n28443 , n14173 );
    xnor g1979 ( n24053 , n25225 , n21867 );
    not g1980 ( n6997 , n3861 );
    not g1981 ( n20017 , n13171 );
    and g1982 ( n16974 , n363 , n16358 );
    and g1983 ( n2123 , n15403 , n16573 );
    xnor g1984 ( n13310 , n20971 , n12607 );
    not g1985 ( n31352 , n17521 );
    and g1986 ( n10801 , n9679 , n4836 );
    and g1987 ( n3038 , n28192 , n7029 );
    xnor g1988 ( n14611 , n15558 , n24464 );
    xor g1989 ( n8401 , n6238 , n19405 );
    or g1990 ( n9408 , n19363 , n8966 );
    not g1991 ( n18484 , n17928 );
    not g1992 ( n466 , n11576 );
    not g1993 ( n2821 , n20231 );
    nor g1994 ( n27447 , n15052 , n29888 );
    not g1995 ( n563 , n20660 );
    and g1996 ( n27340 , n3740 , n23421 );
    or g1997 ( n21608 , n4286 , n10930 );
    not g1998 ( n9002 , n5969 );
    xnor g1999 ( n16146 , n7860 , n20990 );
    and g2000 ( n18616 , n20319 , n11169 );
    xnor g2001 ( n14409 , n746 , n17993 );
    not g2002 ( n18181 , n17024 );
    and g2003 ( n5176 , n12921 , n21519 );
    not g2004 ( n9870 , n16998 );
    not g2005 ( n4155 , n29895 );
    or g2006 ( n9450 , n15172 , n4964 );
    xnor g2007 ( n21842 , n14498 , n8357 );
    or g2008 ( n11024 , n28078 , n7606 );
    or g2009 ( n8343 , n7081 , n27841 );
    and g2010 ( n31947 , n885 , n31291 );
    not g2011 ( n15629 , n17992 );
    buf g2012 ( n20667 , n19770 );
    xnor g2013 ( n10429 , n31591 , n16308 );
    not g2014 ( n24638 , n3131 );
    not g2015 ( n30603 , n5141 );
    or g2016 ( n6618 , n8525 , n15061 );
    xnor g2017 ( n22696 , n22316 , n21466 );
    xnor g2018 ( n20727 , n8554 , n15240 );
    xnor g2019 ( n27951 , n9191 , n29762 );
    or g2020 ( n9429 , n13213 , n27662 );
    and g2021 ( n2184 , n31867 , n29571 );
    not g2022 ( n10400 , n15201 );
    and g2023 ( n23440 , n485 , n17985 );
    xnor g2024 ( n31790 , n5769 , n9845 );
    or g2025 ( n5074 , n17930 , n11313 );
    xnor g2026 ( n16058 , n12764 , n14876 );
    and g2027 ( n26794 , n11905 , n3996 );
    not g2028 ( n8484 , n9831 );
    not g2029 ( n30978 , n6796 );
    and g2030 ( n29594 , n31674 , n25096 );
    or g2031 ( n17128 , n31548 , n20052 );
    and g2032 ( n24263 , n4106 , n15980 );
    nor g2033 ( n22911 , n3062 , n2086 );
    or g2034 ( n12227 , n12453 , n24249 );
    not g2035 ( n8359 , n23417 );
    not g2036 ( n26852 , n21064 );
    or g2037 ( n1673 , n23627 , n8186 );
    not g2038 ( n31255 , n13147 );
    and g2039 ( n773 , n21724 , n12982 );
    and g2040 ( n21437 , n15979 , n9686 );
    and g2041 ( n23356 , n27619 , n29698 );
    not g2042 ( n5191 , n188 );
    and g2043 ( n11516 , n6928 , n7659 );
    xnor g2044 ( n19144 , n13040 , n3949 );
    or g2045 ( n24399 , n1520 , n577 );
    or g2046 ( n23086 , n31129 , n12069 );
    or g2047 ( n13953 , n30052 , n29535 );
    xnor g2048 ( n13270 , n4844 , n24304 );
    or g2049 ( n2927 , n3678 , n27462 );
    not g2050 ( n30572 , n15954 );
    xnor g2051 ( n21170 , n1870 , n13494 );
    not g2052 ( n12899 , n9206 );
    not g2053 ( n22568 , n22809 );
    or g2054 ( n9360 , n9655 , n30601 );
    and g2055 ( n26142 , n18375 , n23768 );
    xnor g2056 ( n11467 , n18253 , n20198 );
    not g2057 ( n25844 , n7611 );
    not g2058 ( n15345 , n1607 );
    xnor g2059 ( n19933 , n3789 , n26117 );
    not g2060 ( n5973 , n13674 );
    xnor g2061 ( n22343 , n28062 , n31837 );
    and g2062 ( n22001 , n6618 , n4770 );
    nor g2063 ( n4386 , n3808 , n23423 );
    or g2064 ( n11818 , n8452 , n463 );
    nor g2065 ( n3853 , n24807 , n8712 );
    not g2066 ( n30130 , n8282 );
    xnor g2067 ( n29693 , n31503 , n22803 );
    not g2068 ( n25170 , n26439 );
    xnor g2069 ( n9390 , n24948 , n19563 );
    or g2070 ( n16834 , n10006 , n20785 );
    or g2071 ( n8193 , n2857 , n21090 );
    xnor g2072 ( n18917 , n4615 , n26408 );
    and g2073 ( n29737 , n14128 , n2346 );
    or g2074 ( n22655 , n7884 , n3544 );
    xnor g2075 ( n15300 , n5110 , n3190 );
    or g2076 ( n18636 , n19226 , n14511 );
    and g2077 ( n21893 , n5077 , n2488 );
    xnor g2078 ( n3877 , n13554 , n10619 );
    xnor g2079 ( n27982 , n21984 , n1218 );
    xnor g2080 ( n10994 , n595 , n134 );
    or g2081 ( n11559 , n3297 , n26601 );
    xnor g2082 ( n11297 , n29128 , n634 );
    or g2083 ( n30451 , n6717 , n24356 );
    xnor g2084 ( n29721 , n16766 , n14161 );
    or g2085 ( n25473 , n3483 , n22997 );
    nor g2086 ( n27814 , n16347 , n12627 );
    and g2087 ( n12366 , n447 , n18948 );
    xnor g2088 ( n30740 , n2372 , n8919 );
    or g2089 ( n14951 , n18305 , n20553 );
    or g2090 ( n20527 , n14280 , n1031 );
    not g2091 ( n22579 , n15711 );
    or g2092 ( n21035 , n9503 , n17456 );
    xor g2093 ( n20020 , n6562 , n22106 );
    or g2094 ( n5119 , n11584 , n29140 );
    xnor g2095 ( n15946 , n2924 , n1980 );
    not g2096 ( n29849 , n27676 );
    or g2097 ( n20124 , n18259 , n6316 );
    or g2098 ( n9648 , n18093 , n10344 );
    and g2099 ( n17690 , n19851 , n5140 );
    xnor g2100 ( n26510 , n2772 , n4845 );
    or g2101 ( n28167 , n19465 , n112 );
    or g2102 ( n13803 , n13770 , n19950 );
    xnor g2103 ( n4402 , n2513 , n16653 );
    nor g2104 ( n15068 , n28417 , n9691 );
    nor g2105 ( n26338 , n13476 , n15818 );
    nor g2106 ( n8959 , n29270 , n4191 );
    not g2107 ( n14267 , n19919 );
    xnor g2108 ( n23156 , n1843 , n15603 );
    xnor g2109 ( n21622 , n11572 , n13359 );
    or g2110 ( n7678 , n8122 , n29787 );
    or g2111 ( n17921 , n26247 , n15635 );
    or g2112 ( n12027 , n25679 , n22954 );
    and g2113 ( n26975 , n17318 , n24122 );
    not g2114 ( n17219 , n20002 );
    xnor g2115 ( n6700 , n1471 , n4249 );
    or g2116 ( n13099 , n4084 , n16903 );
    or g2117 ( n9283 , n22512 , n937 );
    not g2118 ( n22292 , n25492 );
    not g2119 ( n5674 , n9193 );
    and g2120 ( n21693 , n12938 , n20902 );
    not g2121 ( n14159 , n13310 );
    and g2122 ( n8779 , n10436 , n25537 );
    and g2123 ( n1642 , n8181 , n12129 );
    and g2124 ( n8769 , n25706 , n16036 );
    xnor g2125 ( n8760 , n15743 , n4267 );
    or g2126 ( n19588 , n31287 , n10763 );
    xnor g2127 ( n31615 , n31608 , n29747 );
    not g2128 ( n23015 , n31010 );
    nor g2129 ( n22221 , n1232 , n1192 );
    not g2130 ( n24910 , n7241 );
    not g2131 ( n19508 , n20015 );
    nor g2132 ( n3147 , n30649 , n10017 );
    or g2133 ( n27350 , n6267 , n9853 );
    or g2134 ( n16543 , n107 , n16884 );
    nor g2135 ( n16390 , n28856 , n14356 );
    not g2136 ( n4325 , n18275 );
    not g2137 ( n29439 , n29330 );
    not g2138 ( n17330 , n4085 );
    xnor g2139 ( n14668 , n17803 , n9029 );
    xnor g2140 ( n9796 , n6004 , n25428 );
    xor g2141 ( n19797 , n6792 , n17950 );
    not g2142 ( n27004 , n5882 );
    and g2143 ( n3052 , n3397 , n23477 );
    or g2144 ( n30581 , n19511 , n1104 );
    or g2145 ( n26022 , n7110 , n25743 );
    xnor g2146 ( n8387 , n11493 , n14766 );
    or g2147 ( n9433 , n29801 , n26109 );
    and g2148 ( n25128 , n9009 , n30675 );
    or g2149 ( n7436 , n13336 , n23866 );
    and g2150 ( n16897 , n16289 , n1398 );
    nor g2151 ( n7643 , n9973 , n4030 );
    xnor g2152 ( n24563 , n31132 , n12896 );
    xnor g2153 ( n25178 , n30516 , n10786 );
    xnor g2154 ( n2460 , n5638 , n14795 );
    not g2155 ( n4003 , n19549 );
    not g2156 ( n54 , n23639 );
    and g2157 ( n14775 , n28244 , n24726 );
    not g2158 ( n19133 , n1798 );
    or g2159 ( n28660 , n18149 , n19394 );
    xor g2160 ( n17824 , n12295 , n4956 );
    not g2161 ( n12125 , n632 );
    nor g2162 ( n26625 , n25937 , n23504 );
    xnor g2163 ( n23089 , n14950 , n9259 );
    not g2164 ( n911 , n9543 );
    xnor g2165 ( n3880 , n28578 , n12284 );
    xnor g2166 ( n24874 , n18029 , n18644 );
    not g2167 ( n13382 , n3011 );
    and g2168 ( n8866 , n24656 , n19555 );
    nor g2169 ( n4716 , n7345 , n31901 );
    xnor g2170 ( n10037 , n15363 , n20041 );
    or g2171 ( n22740 , n25791 , n19561 );
    and g2172 ( n23566 , n22897 , n17027 );
    or g2173 ( n8658 , n18577 , n26982 );
    not g2174 ( n25832 , n6708 );
    xnor g2175 ( n22460 , n23834 , n13594 );
    or g2176 ( n17275 , n18312 , n19743 );
    or g2177 ( n12089 , n24451 , n18105 );
    not g2178 ( n6951 , n8788 );
    or g2179 ( n13639 , n8938 , n19276 );
    and g2180 ( n30221 , n3985 , n22737 );
    or g2181 ( n28076 , n11881 , n20512 );
    or g2182 ( n15489 , n15952 , n23452 );
    not g2183 ( n26726 , n24416 );
    xnor g2184 ( n18846 , n1192 , n5141 );
    xnor g2185 ( n5757 , n31651 , n7128 );
    not g2186 ( n27005 , n20475 );
    and g2187 ( n16593 , n12291 , n17538 );
    and g2188 ( n14856 , n27032 , n30116 );
    not g2189 ( n16309 , n27513 );
    or g2190 ( n17129 , n25074 , n3528 );
    not g2191 ( n31813 , n14828 );
    and g2192 ( n17481 , n26371 , n20118 );
    not g2193 ( n12980 , n25628 );
    not g2194 ( n31986 , n20708 );
    nor g2195 ( n27505 , n20905 , n28851 );
    not g2196 ( n27585 , n20610 );
    xnor g2197 ( n15998 , n1442 , n14685 );
    xnor g2198 ( n4313 , n15899 , n27566 );
    and g2199 ( n29487 , n6638 , n5548 );
    xnor g2200 ( n14985 , n6522 , n19878 );
    and g2201 ( n16612 , n9648 , n4903 );
    not g2202 ( n18820 , n24522 );
    and g2203 ( n8078 , n134 , n12853 );
    not g2204 ( n29008 , n4570 );
    or g2205 ( n31132 , n2211 , n19469 );
    xnor g2206 ( n16277 , n11929 , n7788 );
    or g2207 ( n30694 , n14446 , n28892 );
    or g2208 ( n2126 , n23642 , n7713 );
    xnor g2209 ( n4659 , n18496 , n7787 );
    xnor g2210 ( n9512 , n13685 , n10114 );
    not g2211 ( n8994 , n793 );
    xnor g2212 ( n4913 , n1039 , n4836 );
    or g2213 ( n7802 , n9835 , n11863 );
    not g2214 ( n10315 , n14992 );
    xnor g2215 ( n16155 , n15646 , n30544 );
    or g2216 ( n2366 , n6733 , n4343 );
    or g2217 ( n20432 , n18766 , n28465 );
    nor g2218 ( n29802 , n5812 , n3677 );
    and g2219 ( n21898 , n10221 , n15956 );
    xor g2220 ( n27236 , n4412 , n30769 );
    not g2221 ( n2462 , n7925 );
    and g2222 ( n19005 , n6966 , n5467 );
    and g2223 ( n31297 , n20191 , n14331 );
    not g2224 ( n15917 , n12783 );
    or g2225 ( n13603 , n6649 , n2992 );
    or g2226 ( n13153 , n31896 , n19569 );
    not g2227 ( n22344 , n3345 );
    or g2228 ( n24656 , n11892 , n28793 );
    xor g2229 ( n27134 , n23454 , n7600 );
    xnor g2230 ( n27772 , n2219 , n6107 );
    xnor g2231 ( n1725 , n22409 , n10377 );
    not g2232 ( n21157 , n7534 );
    xnor g2233 ( n2908 , n23086 , n14305 );
    not g2234 ( n30689 , n20957 );
    and g2235 ( n29367 , n15920 , n4629 );
    xnor g2236 ( n1660 , n9615 , n16402 );
    and g2237 ( n7506 , n20740 , n24944 );
    xnor g2238 ( n616 , n1920 , n21264 );
    or g2239 ( n6812 , n23047 , n7413 );
    xnor g2240 ( n19707 , n31801 , n9849 );
    not g2241 ( n26735 , n2459 );
    or g2242 ( n31670 , n27326 , n24640 );
    not g2243 ( n28381 , n5375 );
    and g2244 ( n30146 , n29223 , n28647 );
    xnor g2245 ( n28625 , n29936 , n4054 );
    or g2246 ( n5053 , n26109 , n29166 );
    and g2247 ( n15585 , n6744 , n7405 );
    or g2248 ( n28692 , n3080 , n2934 );
    not g2249 ( n15531 , n17950 );
    xnor g2250 ( n22182 , n6528 , n26011 );
    and g2251 ( n7121 , n30134 , n191 );
    not g2252 ( n27346 , n259 );
    not g2253 ( n6316 , n2540 );
    xnor g2254 ( n29993 , n23974 , n20145 );
    not g2255 ( n13735 , n10088 );
    xnor g2256 ( n26696 , n27700 , n24561 );
    or g2257 ( n19860 , n29071 , n26117 );
    not g2258 ( n4722 , n27034 );
    xnor g2259 ( n30655 , n29940 , n27046 );
    xnor g2260 ( n30311 , n26255 , n14063 );
    xnor g2261 ( n5270 , n30454 , n14456 );
    not g2262 ( n6849 , n1725 );
    xnor g2263 ( n771 , n20398 , n8017 );
    or g2264 ( n22263 , n12708 , n13882 );
    xnor g2265 ( n26768 , n29882 , n29102 );
    and g2266 ( n23224 , n28730 , n10 );
    or g2267 ( n3351 , n28126 , n4420 );
    not g2268 ( n6936 , n1945 );
    or g2269 ( n29769 , n19995 , n31592 );
    or g2270 ( n12213 , n5436 , n2052 );
    not g2271 ( n26443 , n9476 );
    and g2272 ( n31753 , n13588 , n13500 );
    or g2273 ( n15149 , n21798 , n28539 );
    nor g2274 ( n617 , n11864 , n2449 );
    not g2275 ( n26339 , n26893 );
    xnor g2276 ( n3917 , n19045 , n18224 );
    xnor g2277 ( n9923 , n2063 , n20386 );
    or g2278 ( n22894 , n5770 , n26525 );
    and g2279 ( n11312 , n22812 , n23599 );
    or g2280 ( n27921 , n7624 , n31659 );
    xnor g2281 ( n11839 , n3162 , n30776 );
    xnor g2282 ( n31411 , n19417 , n10304 );
    xnor g2283 ( n15049 , n13626 , n27214 );
    xnor g2284 ( n12867 , n24062 , n2959 );
    not g2285 ( n3727 , n21713 );
    xnor g2286 ( n18510 , n19047 , n29341 );
    and g2287 ( n12068 , n15741 , n16184 );
    or g2288 ( n11356 , n692 , n26101 );
    or g2289 ( n15575 , n31934 , n24700 );
    or g2290 ( n11179 , n22645 , n20611 );
    not g2291 ( n27127 , n29106 );
    not g2292 ( n11475 , n28435 );
    not g2293 ( n5550 , n14955 );
    not g2294 ( n3508 , n21808 );
    not g2295 ( n15427 , n29818 );
    or g2296 ( n14855 , n20232 , n4763 );
    not g2297 ( n27920 , n3396 );
    not g2298 ( n4517 , n5388 );
    and g2299 ( n30235 , n3871 , n26063 );
    not g2300 ( n4489 , n9561 );
    xnor g2301 ( n11255 , n27271 , n13701 );
    nor g2302 ( n29085 , n7414 , n8584 );
    or g2303 ( n9618 , n31179 , n9251 );
    or g2304 ( n26476 , n626 , n15897 );
    xnor g2305 ( n29236 , n24846 , n30704 );
    xnor g2306 ( n19187 , n28797 , n14107 );
    or g2307 ( n24454 , n31357 , n29609 );
    xnor g2308 ( n13674 , n11042 , n29318 );
    xnor g2309 ( n23507 , n14480 , n7017 );
    and g2310 ( n24902 , n20019 , n16675 );
    xnor g2311 ( n31295 , n20217 , n29406 );
    or g2312 ( n3496 , n23440 , n29230 );
    not g2313 ( n1623 , n5801 );
    nor g2314 ( n6959 , n16283 , n24769 );
    not g2315 ( n6104 , n4219 );
    xnor g2316 ( n10055 , n17554 , n11648 );
    xnor g2317 ( n14045 , n1225 , n14712 );
    not g2318 ( n13434 , n21290 );
    xnor g2319 ( n2377 , n24753 , n26603 );
    or g2320 ( n16150 , n24246 , n14376 );
    xnor g2321 ( n3713 , n12418 , n7753 );
    and g2322 ( n14789 , n1050 , n31672 );
    not g2323 ( n5317 , n11788 );
    xnor g2324 ( n9455 , n15691 , n28899 );
    and g2325 ( n28043 , n11732 , n28547 );
    and g2326 ( n17618 , n24791 , n409 );
    not g2327 ( n26627 , n9831 );
    not g2328 ( n24590 , n11495 );
    not g2329 ( n697 , n10883 );
    or g2330 ( n1936 , n16912 , n18887 );
    and g2331 ( n31113 , n20174 , n26955 );
    not g2332 ( n13734 , n15759 );
    or g2333 ( n3918 , n27656 , n1523 );
    and g2334 ( n11436 , n10109 , n30457 );
    xnor g2335 ( n17122 , n15847 , n19356 );
    or g2336 ( n23296 , n1902 , n4457 );
    not g2337 ( n5541 , n4408 );
    not g2338 ( n8796 , n365 );
    and g2339 ( n23535 , n11410 , n31014 );
    or g2340 ( n2923 , n15909 , n77 );
    not g2341 ( n9773 , n29649 );
    nor g2342 ( n25348 , n23126 , n15170 );
    not g2343 ( n17605 , n25091 );
    xnor g2344 ( n7043 , n6190 , n6103 );
    not g2345 ( n11327 , n23019 );
    and g2346 ( n26196 , n13902 , n17305 );
    and g2347 ( n28716 , n10672 , n30914 );
    or g2348 ( n14360 , n8535 , n3537 );
    xnor g2349 ( n24924 , n17176 , n11847 );
    xnor g2350 ( n30590 , n18253 , n16132 );
    or g2351 ( n9761 , n1394 , n11342 );
    and g2352 ( n4363 , n21147 , n13728 );
    xnor g2353 ( n20885 , n445 , n18389 );
    not g2354 ( n28021 , n3119 );
    xor g2355 ( n4960 , n26016 , n6244 );
    not g2356 ( n15238 , n21841 );
    nor g2357 ( n21852 , n26855 , n29061 );
    nor g2358 ( n14306 , n7707 , n12762 );
    or g2359 ( n28345 , n20292 , n23696 );
    not g2360 ( n3085 , n27855 );
    and g2361 ( n21729 , n30284 , n25124 );
    xnor g2362 ( n27157 , n2486 , n17180 );
    or g2363 ( n10011 , n2697 , n7461 );
    or g2364 ( n9558 , n4069 , n28922 );
    and g2365 ( n4549 , n9288 , n28917 );
    not g2366 ( n6364 , n31034 );
    xnor g2367 ( n162 , n30158 , n25242 );
    xnor g2368 ( n20934 , n380 , n10130 );
    xnor g2369 ( n31571 , n7298 , n31433 );
    or g2370 ( n8033 , n13502 , n800 );
    nor g2371 ( n6366 , n5155 , n29971 );
    not g2372 ( n16885 , n28705 );
    or g2373 ( n12512 , n6954 , n29246 );
    nor g2374 ( n17876 , n22512 , n3501 );
    not g2375 ( n797 , n20202 );
    not g2376 ( n18517 , n8004 );
    and g2377 ( n12093 , n12608 , n21630 );
    nor g2378 ( n29433 , n10773 , n17754 );
    or g2379 ( n17769 , n16929 , n5774 );
    not g2380 ( n25195 , n16028 );
    xnor g2381 ( n30903 , n21216 , n30293 );
    and g2382 ( n11888 , n21590 , n27377 );
    or g2383 ( n21103 , n22659 , n16222 );
    and g2384 ( n25044 , n13165 , n23370 );
    and g2385 ( n20087 , n5582 , n3295 );
    and g2386 ( n6193 , n9407 , n6115 );
    xnor g2387 ( n5054 , n5714 , n5254 );
    or g2388 ( n13880 , n651 , n6255 );
    or g2389 ( n28877 , n7758 , n2 );
    and g2390 ( n6389 , n8360 , n29003 );
    nor g2391 ( n6978 , n13616 , n27374 );
    not g2392 ( n10385 , n21535 );
    and g2393 ( n3638 , n502 , n31797 );
    not g2394 ( n4751 , n28864 );
    or g2395 ( n22266 , n14136 , n27242 );
    or g2396 ( n9170 , n18632 , n8257 );
    or g2397 ( n22050 , n21129 , n19519 );
    not g2398 ( n3465 , n25346 );
    xor g2399 ( n17734 , n21581 , n1475 );
    not g2400 ( n8549 , n17085 );
    not g2401 ( n14375 , n11002 );
    not g2402 ( n20633 , n29376 );
    xnor g2403 ( n31990 , n8339 , n19258 );
    or g2404 ( n6625 , n19211 , n7707 );
    not g2405 ( n10979 , n30522 );
    not g2406 ( n9637 , n29349 );
    xnor g2407 ( n7825 , n26510 , n26333 );
    xnor g2408 ( n6902 , n8139 , n14361 );
    nor g2409 ( n11021 , n14390 , n5775 );
    xor g2410 ( n15041 , n6269 , n26765 );
    or g2411 ( n29536 , n9927 , n3497 );
    and g2412 ( n10206 , n10603 , n20475 );
    or g2413 ( n16780 , n24951 , n26017 );
    or g2414 ( n22989 , n10157 , n21886 );
    xnor g2415 ( n30120 , n13600 , n27401 );
    xnor g2416 ( n6403 , n15341 , n9458 );
    xnor g2417 ( n8160 , n21638 , n7351 );
    xor g2418 ( n9788 , n766 , n14323 );
    xnor g2419 ( n1261 , n24388 , n4350 );
    and g2420 ( n21438 , n4976 , n19151 );
    xnor g2421 ( n3482 , n17851 , n891 );
    xnor g2422 ( n16639 , n7934 , n23046 );
    not g2423 ( n28697 , n3080 );
    or g2424 ( n12917 , n26540 , n13088 );
    and g2425 ( n23809 , n1222 , n15859 );
    nor g2426 ( n1988 , n11130 , n15678 );
    not g2427 ( n22260 , n16719 );
    xnor g2428 ( n13041 , n21240 , n18542 );
    not g2429 ( n19633 , n3943 );
    xnor g2430 ( n26998 , n23349 , n21918 );
    xor g2431 ( n945 , n17000 , n25140 );
    or g2432 ( n25086 , n31637 , n8119 );
    not g2433 ( n10005 , n7157 );
    or g2434 ( n16060 , n11446 , n28910 );
    or g2435 ( n19810 , n12312 , n27688 );
    not g2436 ( n8700 , n22256 );
    or g2437 ( n25737 , n24671 , n20372 );
    or g2438 ( n19750 , n2531 , n20103 );
    not g2439 ( n22052 , n1037 );
    or g2440 ( n5461 , n10746 , n29295 );
    xnor g2441 ( n469 , n27222 , n13333 );
    not g2442 ( n17710 , n12634 );
    not g2443 ( n7277 , n763 );
    xnor g2444 ( n5228 , n4847 , n12207 );
    or g2445 ( n25717 , n28777 , n24931 );
    or g2446 ( n790 , n9043 , n26541 );
    not g2447 ( n30071 , n800 );
    nor g2448 ( n27478 , n1980 , n21808 );
    not g2449 ( n4450 , n12131 );
    or g2450 ( n12529 , n19842 , n19688 );
    xnor g2451 ( n9380 , n24392 , n5578 );
    or g2452 ( n19602 , n9472 , n20312 );
    or g2453 ( n25956 , n23561 , n28546 );
    and g2454 ( n17978 , n21811 , n31911 );
    xnor g2455 ( n7070 , n25260 , n16660 );
    or g2456 ( n11637 , n9469 , n22922 );
    or g2457 ( n5157 , n3694 , n2035 );
    and g2458 ( n5422 , n30445 , n30135 );
    xnor g2459 ( n10753 , n1038 , n17550 );
    or g2460 ( n14991 , n4147 , n6673 );
    not g2461 ( n3318 , n26002 );
    nor g2462 ( n14310 , n9282 , n807 );
    and g2463 ( n1598 , n556 , n18332 );
    and g2464 ( n14052 , n16246 , n27879 );
    and g2465 ( n15444 , n13041 , n19366 );
    not g2466 ( n6798 , n6756 );
    not g2467 ( n11950 , n2924 );
    not g2468 ( n26358 , n16873 );
    and g2469 ( n20785 , n20640 , n2161 );
    or g2470 ( n5634 , n28057 , n11499 );
    nor g2471 ( n9456 , n4140 , n170 );
    or g2472 ( n552 , n15411 , n18614 );
    or g2473 ( n29585 , n22432 , n18440 );
    and g2474 ( n21904 , n12250 , n676 );
    nor g2475 ( n5169 , n14391 , n16747 );
    and g2476 ( n30219 , n8037 , n3036 );
    nor g2477 ( n14631 , n11060 , n4174 );
    buf g2478 ( n12979 , n4423 );
    or g2479 ( n25923 , n14477 , n16362 );
    not g2480 ( n19013 , n17801 );
    not g2481 ( n15834 , n19617 );
    and g2482 ( n24864 , n30078 , n2314 );
    xnor g2483 ( n28670 , n15196 , n7938 );
    or g2484 ( n7578 , n16404 , n16583 );
    and g2485 ( n17034 , n691 , n7752 );
    not g2486 ( n27774 , n8773 );
    not g2487 ( n12809 , n28521 );
    nor g2488 ( n341 , n10071 , n10863 );
    xnor g2489 ( n14116 , n23040 , n8834 );
    nor g2490 ( n24599 , n26916 , n4634 );
    nor g2491 ( n19961 , n24394 , n21974 );
    and g2492 ( n29103 , n31605 , n31442 );
    not g2493 ( n27139 , n3567 );
    or g2494 ( n18603 , n29891 , n13393 );
    or g2495 ( n12248 , n19369 , n7116 );
    not g2496 ( n28584 , n10490 );
    nor g2497 ( n1895 , n22867 , n28912 );
    not g2498 ( n29686 , n22141 );
    not g2499 ( n17057 , n14854 );
    xnor g2500 ( n31593 , n3755 , n13604 );
    or g2501 ( n6753 , n5755 , n10390 );
    or g2502 ( n14618 , n3310 , n21859 );
    xnor g2503 ( n10346 , n9271 , n7706 );
    not g2504 ( n8562 , n10842 );
    xnor g2505 ( n8478 , n27926 , n26422 );
    not g2506 ( n7968 , n10488 );
    xnor g2507 ( n21504 , n19538 , n13859 );
    xnor g2508 ( n4127 , n28790 , n16084 );
    xnor g2509 ( n9760 , n28245 , n31092 );
    or g2510 ( n25468 , n28662 , n24057 );
    not g2511 ( n21371 , n21185 );
    not g2512 ( n4299 , n993 );
    not g2513 ( n3540 , n28471 );
    nor g2514 ( n20000 , n28630 , n6327 );
    xnor g2515 ( n3734 , n22122 , n8873 );
    xnor g2516 ( n26255 , n578 , n23532 );
    and g2517 ( n19422 , n27258 , n11375 );
    not g2518 ( n24481 , n13708 );
    not g2519 ( n15536 , n6816 );
    nor g2520 ( n10941 , n13221 , n24944 );
    or g2521 ( n19639 , n30371 , n18044 );
    not g2522 ( n21257 , n14197 );
    or g2523 ( n1506 , n29521 , n21698 );
    not g2524 ( n9766 , n3668 );
    not g2525 ( n27454 , n31546 );
    or g2526 ( n7635 , n180 , n15065 );
    xnor g2527 ( n30829 , n20816 , n17802 );
    xnor g2528 ( n20088 , n15342 , n17457 );
    or g2529 ( n7699 , n14534 , n14839 );
    nor g2530 ( n24055 , n14555 , n15648 );
    xnor g2531 ( n25251 , n27956 , n9273 );
    xnor g2532 ( n15924 , n775 , n30287 );
    or g2533 ( n12302 , n30300 , n21171 );
    xnor g2534 ( n16853 , n2792 , n11357 );
    and g2535 ( n29696 , n17139 , n14727 );
    xnor g2536 ( n15780 , n5243 , n29836 );
    or g2537 ( n23747 , n4572 , n7121 );
    not g2538 ( n8111 , n11197 );
    not g2539 ( n2311 , n17149 );
    xnor g2540 ( n4774 , n10406 , n18977 );
    or g2541 ( n23421 , n26004 , n2324 );
    and g2542 ( n20734 , n18962 , n10517 );
    xor g2543 ( n1147 , n22245 , n2466 );
    and g2544 ( n11184 , n455 , n26608 );
    and g2545 ( n16769 , n2132 , n7501 );
    xnor g2546 ( n23613 , n29656 , n13054 );
    and g2547 ( n6221 , n14543 , n28091 );
    and g2548 ( n11426 , n4456 , n17837 );
    xnor g2549 ( n8251 , n22484 , n13546 );
    xnor g2550 ( n18395 , n17399 , n5448 );
    or g2551 ( n6588 , n29764 , n2315 );
    or g2552 ( n30826 , n29878 , n9096 );
    or g2553 ( n19551 , n25422 , n606 );
    xnor g2554 ( n14741 , n21066 , n26178 );
    not g2555 ( n19937 , n23679 );
    xnor g2556 ( n31390 , n26618 , n31456 );
    or g2557 ( n26014 , n11054 , n28484 );
    not g2558 ( n21252 , n6500 );
    and g2559 ( n24713 , n7041 , n31507 );
    xnor g2560 ( n16775 , n23447 , n1062 );
    and g2561 ( n11522 , n28113 , n14949 );
    nor g2562 ( n10036 , n24712 , n835 );
    buf g2563 ( n7068 , n22216 );
    and g2564 ( n4986 , n27047 , n8658 );
    or g2565 ( n8889 , n10057 , n21077 );
    and g2566 ( n22459 , n22191 , n20816 );
    not g2567 ( n28413 , n7904 );
    not g2568 ( n22650 , n265 );
    or g2569 ( n25181 , n28328 , n30673 );
    and g2570 ( n27083 , n31814 , n13931 );
    and g2571 ( n8855 , n28436 , n22137 );
    or g2572 ( n16905 , n27951 , n17102 );
    or g2573 ( n13331 , n26115 , n21960 );
    not g2574 ( n2219 , n26795 );
    xnor g2575 ( n9526 , n10096 , n28936 );
    not g2576 ( n10810 , n19566 );
    not g2577 ( n21476 , n8415 );
    xnor g2578 ( n21156 , n31044 , n7392 );
    xnor g2579 ( n21067 , n29349 , n5773 );
    or g2580 ( n14258 , n19382 , n2695 );
    or g2581 ( n16681 , n5029 , n17243 );
    and g2582 ( n6212 , n11313 , n22300 );
    not g2583 ( n1668 , n14477 );
    or g2584 ( n15404 , n4119 , n4261 );
    not g2585 ( n23725 , n20825 );
    xnor g2586 ( n22369 , n25216 , n24482 );
    xnor g2587 ( n28787 , n16553 , n3221 );
    not g2588 ( n10851 , n19924 );
    or g2589 ( n16138 , n14782 , n2121 );
    or g2590 ( n8740 , n22326 , n23103 );
    nor g2591 ( n19751 , n26748 , n25481 );
    xnor g2592 ( n31822 , n4010 , n4504 );
    or g2593 ( n25767 , n682 , n9764 );
    xor g2594 ( n3189 , n23897 , n9843 );
    nor g2595 ( n31490 , n18349 , n8678 );
    and g2596 ( n13128 , n8777 , n27496 );
    or g2597 ( n13072 , n1776 , n26587 );
    or g2598 ( n24475 , n30677 , n7337 );
    and g2599 ( n1389 , n11320 , n250 );
    not g2600 ( n16791 , n31178 );
    and g2601 ( n22150 , n5124 , n18799 );
    or g2602 ( n8135 , n19319 , n12144 );
    or g2603 ( n11532 , n12526 , n22915 );
    xnor g2604 ( n6889 , n24443 , n5077 );
    or g2605 ( n3317 , n14670 , n11576 );
    xnor g2606 ( n17801 , n24393 , n14257 );
    nor g2607 ( n13746 , n31503 , n18421 );
    xnor g2608 ( n26955 , n8441 , n9111 );
    or g2609 ( n7579 , n1331 , n6365 );
    not g2610 ( n1508 , n4751 );
    not g2611 ( n10249 , n22778 );
    or g2612 ( n1905 , n28070 , n7298 );
    xnor g2613 ( n22726 , n19160 , n3056 );
    not g2614 ( n17557 , n21010 );
    not g2615 ( n26087 , n22832 );
    nor g2616 ( n29768 , n9574 , n31013 );
    nor g2617 ( n4557 , n28081 , n3004 );
    and g2618 ( n2440 , n7327 , n17083 );
    nor g2619 ( n3168 , n7757 , n10712 );
    or g2620 ( n19115 , n30900 , n20921 );
    and g2621 ( n22480 , n20658 , n10279 );
    or g2622 ( n10611 , n22269 , n13250 );
    not g2623 ( n16928 , n7534 );
    xnor g2624 ( n23284 , n9720 , n2231 );
    not g2625 ( n1643 , n27 );
    and g2626 ( n17777 , n9678 , n23005 );
    and g2627 ( n11256 , n31383 , n3629 );
    xnor g2628 ( n4516 , n16256 , n28507 );
    xnor g2629 ( n9945 , n23953 , n29611 );
    or g2630 ( n25038 , n28525 , n9701 );
    and g2631 ( n21328 , n4639 , n10178 );
    and g2632 ( n16443 , n5194 , n29119 );
    or g2633 ( n14810 , n3077 , n5917 );
    or g2634 ( n29300 , n25442 , n10660 );
    or g2635 ( n20979 , n11462 , n2862 );
    or g2636 ( n11638 , n2963 , n24459 );
    not g2637 ( n17343 , n17480 );
    not g2638 ( n13356 , n17448 );
    not g2639 ( n28022 , n30326 );
    nor g2640 ( n22539 , n8677 , n10970 );
    xnor g2641 ( n11098 , n23680 , n4349 );
    not g2642 ( n192 , n2259 );
    not g2643 ( n28453 , n10433 );
    and g2644 ( n6421 , n25762 , n6774 );
    xnor g2645 ( n30679 , n12852 , n3248 );
    or g2646 ( n23367 , n11018 , n3146 );
    xnor g2647 ( n8999 , n5353 , n1122 );
    or g2648 ( n10983 , n7034 , n14460 );
    nor g2649 ( n16527 , n9044 , n31644 );
    or g2650 ( n10604 , n28904 , n29975 );
    xnor g2651 ( n16270 , n20156 , n23138 );
    or g2652 ( n26463 , n11991 , n13024 );
    not g2653 ( n30853 , n11323 );
    xor g2654 ( n7343 , n8112 , n13152 );
    and g2655 ( n22109 , n6015 , n29529 );
    or g2656 ( n11003 , n22845 , n27362 );
    or g2657 ( n6829 , n28388 , n16325 );
    not g2658 ( n29659 , n1497 );
    not g2659 ( n15064 , n24598 );
    or g2660 ( n13567 , n27375 , n27858 );
    not g2661 ( n27761 , n21372 );
    and g2662 ( n13882 , n17404 , n25501 );
    xnor g2663 ( n5655 , n1916 , n19584 );
    not g2664 ( n24014 , n15127 );
    xnor g2665 ( n10723 , n16740 , n21869 );
    or g2666 ( n14232 , n304 , n23442 );
    and g2667 ( n20396 , n17878 , n15342 );
    xnor g2668 ( n24586 , n3238 , n11370 );
    not g2669 ( n26902 , n21070 );
    not g2670 ( n11677 , n19549 );
    or g2671 ( n17627 , n2554 , n2029 );
    or g2672 ( n19266 , n445 , n5150 );
    or g2673 ( n5947 , n190 , n11148 );
    not g2674 ( n11957 , n29855 );
    buf g2675 ( n5113 , n14630 );
    xnor g2676 ( n28858 , n2201 , n17103 );
    nor g2677 ( n22991 , n12293 , n21919 );
    not g2678 ( n4918 , n10562 );
    or g2679 ( n28916 , n7630 , n2742 );
    xnor g2680 ( n13480 , n25157 , n10196 );
    not g2681 ( n7496 , n26052 );
    not g2682 ( n6921 , n15915 );
    xnor g2683 ( n29126 , n31108 , n29615 );
    xnor g2684 ( n27506 , n19623 , n13812 );
    buf g2685 ( n24630 , n17530 );
    and g2686 ( n31522 , n1890 , n29843 );
    or g2687 ( n207 , n28301 , n24341 );
    not g2688 ( n12282 , n8063 );
    xnor g2689 ( n31181 , n8169 , n4403 );
    not g2690 ( n21881 , n4813 );
    xnor g2691 ( n5736 , n852 , n19655 );
    not g2692 ( n2182 , n3794 );
    xnor g2693 ( n3202 , n8138 , n15835 );
    or g2694 ( n10894 , n25889 , n5881 );
    not g2695 ( n20854 , n31896 );
    or g2696 ( n3989 , n14377 , n10514 );
    and g2697 ( n1356 , n29453 , n19158 );
    not g2698 ( n20283 , n9925 );
    not g2699 ( n9533 , n30287 );
    nor g2700 ( n26484 , n14119 , n7563 );
    and g2701 ( n1248 , n21907 , n630 );
    xnor g2702 ( n16893 , n19296 , n18107 );
    xnor g2703 ( n22342 , n6236 , n2753 );
    xnor g2704 ( n8365 , n20477 , n799 );
    not g2705 ( n21696 , n17124 );
    or g2706 ( n19653 , n18317 , n16874 );
    xnor g2707 ( n8393 , n19790 , n24988 );
    not g2708 ( n24583 , n9616 );
    xnor g2709 ( n21895 , n21122 , n7655 );
    not g2710 ( n22163 , n12953 );
    not g2711 ( n14915 , n11932 );
    xnor g2712 ( n24036 , n27064 , n8873 );
    or g2713 ( n3756 , n16731 , n4189 );
    and g2714 ( n16666 , n3389 , n13972 );
    xnor g2715 ( n213 , n12051 , n14121 );
    or g2716 ( n5553 , n20178 , n23142 );
    or g2717 ( n26516 , n15010 , n3991 );
    not g2718 ( n29888 , n3955 );
    nor g2719 ( n17353 , n11906 , n13482 );
    xnor g2720 ( n5999 , n31773 , n3907 );
    xnor g2721 ( n28145 , n556 , n2061 );
    and g2722 ( n2859 , n28560 , n26556 );
    not g2723 ( n23428 , n14221 );
    not g2724 ( n20994 , n11800 );
    and g2725 ( n12104 , n6474 , n3501 );
    nor g2726 ( n8716 , n25980 , n25558 );
    not g2727 ( n10805 , n13162 );
    and g2728 ( n25782 , n12461 , n12854 );
    and g2729 ( n14959 , n12893 , n10748 );
    or g2730 ( n9268 , n16650 , n17012 );
    and g2731 ( n31778 , n5079 , n17426 );
    xnor g2732 ( n20171 , n2415 , n8699 );
    nor g2733 ( n4788 , n22114 , n8852 );
    not g2734 ( n21496 , n17906 );
    nor g2735 ( n26009 , n13554 , n11737 );
    xor g2736 ( n8143 , n23103 , n10624 );
    buf g2737 ( n28712 , n22358 );
    and g2738 ( n4818 , n30975 , n2849 );
    or g2739 ( n11942 , n30593 , n10129 );
    or g2740 ( n17939 , n12920 , n15081 );
    and g2741 ( n615 , n12341 , n6609 );
    not g2742 ( n6438 , n7922 );
    not g2743 ( n704 , n14836 );
    or g2744 ( n8325 , n14552 , n14551 );
    xnor g2745 ( n24717 , n8986 , n31889 );
    xnor g2746 ( n16661 , n8351 , n28599 );
    and g2747 ( n11883 , n18395 , n28445 );
    xnor g2748 ( n20279 , n17360 , n11128 );
    and g2749 ( n13890 , n1947 , n29325 );
    or g2750 ( n29344 , n11413 , n28069 );
    or g2751 ( n29551 , n20465 , n7941 );
    not g2752 ( n291 , n20040 );
    or g2753 ( n26361 , n10979 , n772 );
    xnor g2754 ( n11338 , n11481 , n31376 );
    and g2755 ( n2066 , n7074 , n20661 );
    not g2756 ( n24792 , n30323 );
    xnor g2757 ( n1811 , n27747 , n29816 );
    or g2758 ( n10535 , n11368 , n28767 );
    not g2759 ( n4102 , n19036 );
    xor g2760 ( n12660 , n8745 , n14011 );
    nor g2761 ( n8504 , n25031 , n14403 );
    not g2762 ( n19783 , n31214 );
    not g2763 ( n8411 , n21777 );
    not g2764 ( n21996 , n21547 );
    and g2765 ( n19171 , n7244 , n8363 );
    not g2766 ( n21394 , n5417 );
    or g2767 ( n11229 , n3349 , n4071 );
    or g2768 ( n19377 , n11855 , n19454 );
    and g2769 ( n29115 , n4461 , n13884 );
    nor g2770 ( n7630 , n7434 , n22512 );
    and g2771 ( n20606 , n15653 , n4314 );
    not g2772 ( n1903 , n17832 );
    or g2773 ( n711 , n5660 , n26183 );
    or g2774 ( n14531 , n5351 , n20007 );
    not g2775 ( n23355 , n13859 );
    nor g2776 ( n25932 , n22235 , n27359 );
    xnor g2777 ( n3906 , n22984 , n10498 );
    nor g2778 ( n1478 , n29830 , n15132 );
    nor g2779 ( n30487 , n6667 , n2984 );
    nor g2780 ( n28484 , n12384 , n4706 );
    and g2781 ( n20605 , n27353 , n29722 );
    xnor g2782 ( n9909 , n21318 , n7113 );
    not g2783 ( n3068 , n1137 );
    xnor g2784 ( n3369 , n29871 , n5313 );
    and g2785 ( n16993 , n16423 , n1436 );
    and g2786 ( n4759 , n2238 , n4428 );
    and g2787 ( n18466 , n1666 , n7206 );
    or g2788 ( n5980 , n3216 , n22872 );
    xnor g2789 ( n29528 , n20823 , n20453 );
    xnor g2790 ( n16384 , n22629 , n30477 );
    xnor g2791 ( n21177 , n9767 , n10288 );
    or g2792 ( n31022 , n11849 , n8877 );
    or g2793 ( n9539 , n15232 , n12971 );
    not g2794 ( n31923 , n2728 );
    not g2795 ( n22326 , n19004 );
    xnor g2796 ( n19452 , n13623 , n21622 );
    buf g2797 ( n8705 , n15162 );
    and g2798 ( n28751 , n436 , n26360 );
    and g2799 ( n31434 , n7097 , n26132 );
    or g2800 ( n1496 , n8834 , n6123 );
    or g2801 ( n17810 , n28974 , n7649 );
    xnor g2802 ( n13940 , n3765 , n10158 );
    not g2803 ( n26323 , n15838 );
    and g2804 ( n5173 , n27194 , n14891 );
    and g2805 ( n8437 , n9112 , n8102 );
    and g2806 ( n10257 , n31930 , n25276 );
    not g2807 ( n22657 , n17595 );
    xnor g2808 ( n14601 , n12984 , n23582 );
    not g2809 ( n25087 , n29994 );
    xnor g2810 ( n8414 , n12999 , n4568 );
    or g2811 ( n16503 , n18677 , n15189 );
    and g2812 ( n28819 , n7635 , n24654 );
    or g2813 ( n5291 , n14159 , n2751 );
    or g2814 ( n9090 , n25972 , n23060 );
    nor g2815 ( n13720 , n24369 , n15836 );
    xnor g2816 ( n6645 , n10108 , n30505 );
    not g2817 ( n13998 , n12946 );
    not g2818 ( n10378 , n3310 );
    not g2819 ( n27715 , n9619 );
    or g2820 ( n20127 , n5788 , n22595 );
    xnor g2821 ( n25310 , n32026 , n10072 );
    not g2822 ( n23780 , n13470 );
    xnor g2823 ( n29308 , n3636 , n16387 );
    not g2824 ( n6435 , n20519 );
    not g2825 ( n4268 , n23673 );
    xnor g2826 ( n10145 , n31174 , n12689 );
    or g2827 ( n29092 , n28180 , n19105 );
    and g2828 ( n6044 , n3269 , n4196 );
    or g2829 ( n14973 , n6222 , n22557 );
    or g2830 ( n30855 , n8264 , n16736 );
    not g2831 ( n28201 , n12233 );
    not g2832 ( n27135 , n24512 );
    not g2833 ( n6969 , n25995 );
    or g2834 ( n26311 , n1277 , n17222 );
    xnor g2835 ( n17568 , n23017 , n10619 );
    xnor g2836 ( n290 , n2139 , n29351 );
    or g2837 ( n14756 , n11487 , n10540 );
    xnor g2838 ( n4625 , n29535 , n4288 );
    xnor g2839 ( n4468 , n6524 , n27839 );
    xnor g2840 ( n4374 , n16388 , n27714 );
    or g2841 ( n31690 , n16301 , n5343 );
    nor g2842 ( n24368 , n28419 , n6359 );
    nor g2843 ( n17320 , n10001 , n29474 );
    not g2844 ( n2509 , n23957 );
    and g2845 ( n4430 , n2418 , n8218 );
    not g2846 ( n3747 , n27681 );
    or g2847 ( n2489 , n18203 , n24858 );
    or g2848 ( n16067 , n10331 , n27644 );
    xnor g2849 ( n25917 , n5234 , n15782 );
    xnor g2850 ( n28338 , n19445 , n29818 );
    xnor g2851 ( n17847 , n4723 , n7867 );
    and g2852 ( n4687 , n24225 , n2528 );
    or g2853 ( n31272 , n11863 , n23725 );
    not g2854 ( n31635 , n3932 );
    xor g2855 ( n16448 , n12093 , n21017 );
    or g2856 ( n10821 , n6807 , n11819 );
    or g2857 ( n3555 , n8885 , n12228 );
    nor g2858 ( n5365 , n25585 , n25976 );
    or g2859 ( n27584 , n22323 , n25471 );
    xnor g2860 ( n14945 , n1616 , n9835 );
    nor g2861 ( n13109 , n2818 , n9758 );
    nor g2862 ( n22900 , n908 , n31211 );
    and g2863 ( n14299 , n20133 , n14181 );
    or g2864 ( n12864 , n29106 , n1550 );
    or g2865 ( n19147 , n3398 , n26366 );
    and g2866 ( n24519 , n14653 , n30229 );
    xnor g2867 ( n10736 , n25897 , n2809 );
    xnor g2868 ( n14300 , n25051 , n17166 );
    not g2869 ( n15243 , n18989 );
    and g2870 ( n24636 , n14978 , n3072 );
    and g2871 ( n28585 , n19697 , n1071 );
    not g2872 ( n31417 , n25543 );
    xnor g2873 ( n14989 , n7725 , n29693 );
    and g2874 ( n8459 , n13639 , n14247 );
    nor g2875 ( n29029 , n31591 , n16308 );
    not g2876 ( n30046 , n10474 );
    or g2877 ( n25030 , n19673 , n5413 );
    or g2878 ( n1034 , n26393 , n581 );
    not g2879 ( n28210 , n18992 );
    xnor g2880 ( n21286 , n21309 , n15744 );
    xnor g2881 ( n31421 , n25101 , n4396 );
    and g2882 ( n26910 , n16583 , n29069 );
    xor g2883 ( n29908 , n31355 , n3614 );
    or g2884 ( n18799 , n8586 , n5822 );
    not g2885 ( n24951 , n26689 );
    or g2886 ( n18826 , n7314 , n30254 );
    not g2887 ( n12241 , n10871 );
    and g2888 ( n30483 , n18226 , n19866 );
    and g2889 ( n29479 , n28897 , n20259 );
    or g2890 ( n7756 , n14769 , n17949 );
    or g2891 ( n25623 , n29615 , n29990 );
    nor g2892 ( n20949 , n26886 , n8821 );
    xnor g2893 ( n6498 , n15010 , n11060 );
    not g2894 ( n23437 , n18253 );
    not g2895 ( n2520 , n24016 );
    not g2896 ( n20227 , n1368 );
    not g2897 ( n26486 , n28763 );
    or g2898 ( n16515 , n24852 , n14623 );
    not g2899 ( n1363 , n27544 );
    not g2900 ( n8246 , n4901 );
    or g2901 ( n7840 , n29384 , n28325 );
    and g2902 ( n2931 , n14578 , n21419 );
    nor g2903 ( n8547 , n5361 , n8931 );
    not g2904 ( n8195 , n25330 );
    not g2905 ( n21661 , n8940 );
    and g2906 ( n25032 , n11852 , n28828 );
    xnor g2907 ( n16551 , n26901 , n21464 );
    not g2908 ( n31416 , n24138 );
    or g2909 ( n8511 , n11155 , n1058 );
    or g2910 ( n17958 , n31439 , n20899 );
    not g2911 ( n6629 , n23490 );
    nor g2912 ( n7356 , n21708 , n12241 );
    xnor g2913 ( n2577 , n1482 , n12507 );
    xnor g2914 ( n24851 , n20327 , n14160 );
    not g2915 ( n16139 , n5262 );
    or g2916 ( n4693 , n17220 , n19590 );
    or g2917 ( n3128 , n22250 , n7415 );
    not g2918 ( n840 , n14821 );
    xnor g2919 ( n25968 , n26509 , n14774 );
    not g2920 ( n8678 , n13233 );
    xnor g2921 ( n13871 , n24696 , n14438 );
    not g2922 ( n18550 , n5110 );
    xnor g2923 ( n10455 , n15189 , n25156 );
    or g2924 ( n10976 , n5545 , n28551 );
    not g2925 ( n7549 , n27401 );
    nor g2926 ( n15655 , n24446 , n9446 );
    not g2927 ( n5744 , n29000 );
    and g2928 ( n8965 , n15559 , n20041 );
    xnor g2929 ( n1964 , n29132 , n28634 );
    and g2930 ( n12693 , n1852 , n31929 );
    xnor g2931 ( n15797 , n31005 , n16438 );
    and g2932 ( n9366 , n13030 , n13823 );
    and g2933 ( n16480 , n15985 , n9089 );
    and g2934 ( n11625 , n29523 , n18433 );
    or g2935 ( n2427 , n23023 , n6340 );
    not g2936 ( n2122 , n24909 );
    nor g2937 ( n25163 , n11795 , n17200 );
    xnor g2938 ( n10299 , n29793 , n26072 );
    and g2939 ( n4 , n5053 , n4369 );
    not g2940 ( n24081 , n12012 );
    xnor g2941 ( n3196 , n18450 , n346 );
    and g2942 ( n28868 , n11525 , n5123 );
    xnor g2943 ( n1565 , n24 , n21186 );
    nor g2944 ( n12574 , n8457 , n3067 );
    not g2945 ( n11899 , n22922 );
    not g2946 ( n13317 , n567 );
    or g2947 ( n10798 , n2346 , n10241 );
    nor g2948 ( n11092 , n10673 , n5114 );
    not g2949 ( n12892 , n3213 );
    and g2950 ( n9357 , n7013 , n655 );
    xnor g2951 ( n20595 , n12945 , n1602 );
    xnor g2952 ( n27836 , n23823 , n20442 );
    xnor g2953 ( n4422 , n20731 , n28975 );
    xnor g2954 ( n11526 , n8855 , n26251 );
    or g2955 ( n11463 , n13703 , n19646 );
    and g2956 ( n24495 , n3945 , n19066 );
    xnor g2957 ( n16950 , n7495 , n20155 );
    xnor g2958 ( n28626 , n28976 , n4409 );
    or g2959 ( n12844 , n11663 , n12857 );
    and g2960 ( n148 , n15874 , n8629 );
    nor g2961 ( n521 , n19405 , n14513 );
    or g2962 ( n3470 , n25699 , n12479 );
    xnor g2963 ( n17174 , n21603 , n30936 );
    or g2964 ( n4726 , n30569 , n6187 );
    or g2965 ( n26086 , n26909 , n29915 );
    or g2966 ( n27887 , n23305 , n2063 );
    or g2967 ( n7832 , n13983 , n18259 );
    or g2968 ( n16992 , n6534 , n19594 );
    not g2969 ( n6783 , n18509 );
    and g2970 ( n13523 , n5051 , n7521 );
    not g2971 ( n7563 , n14601 );
    xnor g2972 ( n11293 , n24939 , n19538 );
    xnor g2973 ( n30236 , n24163 , n906 );
    not g2974 ( n19566 , n27842 );
    or g2975 ( n20852 , n6132 , n4896 );
    or g2976 ( n20685 , n10034 , n1100 );
    xnor g2977 ( n29792 , n12444 , n26376 );
    nor g2978 ( n2573 , n21310 , n15361 );
    or g2979 ( n15239 , n286 , n31472 );
    and g2980 ( n25390 , n20651 , n9074 );
    not g2981 ( n24594 , n24926 );
    xnor g2982 ( n18479 , n1969 , n30667 );
    not g2983 ( n3911 , n31915 );
    or g2984 ( n28619 , n24377 , n26853 );
    xnor g2985 ( n14160 , n22275 , n20337 );
    not g2986 ( n13241 , n12781 );
    or g2987 ( n2345 , n19696 , n28232 );
    xnor g2988 ( n19680 , n8655 , n17368 );
    or g2989 ( n30292 , n12055 , n29507 );
    xnor g2990 ( n27011 , n4759 , n20390 );
    or g2991 ( n24176 , n6780 , n11595 );
    or g2992 ( n1789 , n19039 , n14706 );
    not g2993 ( n5545 , n30090 );
    or g2994 ( n9982 , n23842 , n17743 );
    not g2995 ( n20543 , n1311 );
    or g2996 ( n7614 , n12859 , n14082 );
    or g2997 ( n13787 , n3767 , n2557 );
    not g2998 ( n17221 , n27962 );
    not g2999 ( n16436 , n18087 );
    not g3000 ( n31318 , n13111 );
    or g3001 ( n539 , n19628 , n354 );
    or g3002 ( n5894 , n28427 , n29879 );
    and g3003 ( n17369 , n11875 , n14293 );
    not g3004 ( n15651 , n1020 );
    or g3005 ( n20189 , n29108 , n28390 );
    xnor g3006 ( n8596 , n18856 , n6940 );
    not g3007 ( n27952 , n31702 );
    or g3008 ( n27808 , n19957 , n9256 );
    xnor g3009 ( n8922 , n13957 , n15342 );
    or g3010 ( n11454 , n27686 , n12532 );
    or g3011 ( n1843 , n2338 , n1658 );
    or g3012 ( n14404 , n31258 , n1531 );
    not g3013 ( n6374 , n21104 );
    not g3014 ( n6533 , n23189 );
    and g3015 ( n1641 , n17967 , n27328 );
    not g3016 ( n12014 , n12998 );
    not g3017 ( n21719 , n3013 );
    nor g3018 ( n8147 , n9021 , n23285 );
    not g3019 ( n28919 , n22748 );
    xnor g3020 ( n1701 , n12398 , n14035 );
    or g3021 ( n8115 , n9744 , n17506 );
    xnor g3022 ( n25428 , n3959 , n5938 );
    not g3023 ( n13328 , n17051 );
    not g3024 ( n30187 , n5062 );
    or g3025 ( n28927 , n13762 , n14771 );
    or g3026 ( n21361 , n6527 , n10600 );
    xnor g3027 ( n1312 , n16936 , n29434 );
    not g3028 ( n26756 , n8782 );
    xnor g3029 ( n15231 , n23553 , n30474 );
    xnor g3030 ( n17249 , n29965 , n26620 );
    xnor g3031 ( n4745 , n24410 , n22849 );
    xnor g3032 ( n4131 , n17585 , n20486 );
    or g3033 ( n14442 , n603 , n26112 );
    or g3034 ( n29231 , n31601 , n21434 );
    and g3035 ( n14349 , n27392 , n3768 );
    xnor g3036 ( n13453 , n31569 , n10971 );
    xnor g3037 ( n31948 , n28856 , n14356 );
    or g3038 ( n24458 , n18807 , n18053 );
    and g3039 ( n18280 , n11605 , n27908 );
    xnor g3040 ( n15336 , n27682 , n9782 );
    not g3041 ( n2261 , n28109 );
    and g3042 ( n4574 , n3122 , n23109 );
    xnor g3043 ( n18701 , n17745 , n12920 );
    or g3044 ( n10099 , n25479 , n22562 );
    buf g3045 ( n5561 , n734 );
    not g3046 ( n2308 , n23410 );
    xnor g3047 ( n5640 , n23432 , n492 );
    xnor g3048 ( n15380 , n19432 , n11232 );
    and g3049 ( n14295 , n10345 , n5344 );
    not g3050 ( n25176 , n24056 );
    not g3051 ( n19103 , n17786 );
    or g3052 ( n630 , n1632 , n12912 );
    or g3053 ( n6640 , n12744 , n16480 );
    xor g3054 ( n13136 , n14312 , n19251 );
    and g3055 ( n8717 , n30615 , n10162 );
    not g3056 ( n29091 , n14761 );
    and g3057 ( n30533 , n31592 , n19995 );
    or g3058 ( n663 , n29600 , n10560 );
    or g3059 ( n29087 , n21466 , n14379 );
    or g3060 ( n7036 , n16692 , n18660 );
    and g3061 ( n20529 , n12668 , n29471 );
    xnor g3062 ( n6729 , n6182 , n25415 );
    not g3063 ( n9792 , n23092 );
    xnor g3064 ( n14095 , n14035 , n154 );
    nor g3065 ( n2754 , n12242 , n9509 );
    or g3066 ( n10149 , n25868 , n29685 );
    xnor g3067 ( n10229 , n20930 , n20185 );
    not g3068 ( n26294 , n19619 );
    or g3069 ( n18923 , n28087 , n19492 );
    not g3070 ( n11795 , n22075 );
    xnor g3071 ( n15421 , n20655 , n24909 );
    xnor g3072 ( n17374 , n26444 , n26834 );
    or g3073 ( n24347 , n21181 , n26818 );
    and g3074 ( n2409 , n26499 , n11086 );
    or g3075 ( n12110 , n31606 , n30990 );
    nor g3076 ( n25633 , n4559 , n15057 );
    not g3077 ( n13110 , n12747 );
    nor g3078 ( n11034 , n12072 , n8897 );
    or g3079 ( n6499 , n10253 , n22480 );
    nor g3080 ( n733 , n18078 , n30992 );
    or g3081 ( n18032 , n21786 , n475 );
    xnor g3082 ( n23858 , n14447 , n20815 );
    and g3083 ( n14103 , n23424 , n15473 );
    or g3084 ( n7816 , n15342 , n11624 );
    and g3085 ( n25402 , n31125 , n11325 );
    not g3086 ( n22858 , n9604 );
    not g3087 ( n24917 , n29447 );
    not g3088 ( n30756 , n7525 );
    not g3089 ( n31009 , n30245 );
    or g3090 ( n15902 , n6024 , n16677 );
    xnor g3091 ( n24255 , n11240 , n6833 );
    or g3092 ( n19697 , n25297 , n16875 );
    or g3093 ( n868 , n3036 , n11573 );
    and g3094 ( n12889 , n31276 , n19010 );
    or g3095 ( n10420 , n18587 , n1860 );
    xnor g3096 ( n3478 , n13247 , n9486 );
    not g3097 ( n27343 , n12312 );
    not g3098 ( n30497 , n30717 );
    and g3099 ( n6134 , n6886 , n2281 );
    or g3100 ( n8248 , n23934 , n1232 );
    or g3101 ( n13245 , n4255 , n18657 );
    not g3102 ( n11112 , n24290 );
    xnor g3103 ( n26505 , n20134 , n25407 );
    or g3104 ( n723 , n9209 , n12370 );
    xnor g3105 ( n16306 , n10025 , n12090 );
    or g3106 ( n30217 , n24657 , n10695 );
    or g3107 ( n11087 , n25902 , n26657 );
    or g3108 ( n27426 , n12743 , n17205 );
    or g3109 ( n31971 , n30211 , n958 );
    xnor g3110 ( n17065 , n23023 , n26700 );
    or g3111 ( n9748 , n12784 , n16271 );
    not g3112 ( n30554 , n28588 );
    nor g3113 ( n15966 , n12999 , n23505 );
    not g3114 ( n28203 , n15849 );
    not g3115 ( n23253 , n3664 );
    or g3116 ( n29328 , n81 , n19535 );
    or g3117 ( n7712 , n4653 , n24563 );
    nor g3118 ( n355 , n14527 , n14338 );
    xnor g3119 ( n8368 , n27363 , n11467 );
    or g3120 ( n3226 , n5367 , n11334 );
    xnor g3121 ( n7990 , n30310 , n29418 );
    nor g3122 ( n7287 , n16583 , n13061 );
    and g3123 ( n27052 , n9056 , n14003 );
    xnor g3124 ( n22237 , n19046 , n591 );
    xnor g3125 ( n6103 , n25388 , n30414 );
    or g3126 ( n18835 , n610 , n11741 );
    not g3127 ( n17750 , n30568 );
    xnor g3128 ( n17814 , n9473 , n18678 );
    xnor g3129 ( n28298 , n31036 , n7243 );
    or g3130 ( n2495 , n13936 , n12022 );
    xnor g3131 ( n28849 , n26254 , n12426 );
    xnor g3132 ( n18413 , n10900 , n26565 );
    xor g3133 ( n1575 , n26316 , n11771 );
    not g3134 ( n16161 , n19339 );
    xnor g3135 ( n30711 , n21948 , n6169 );
    xnor g3136 ( n18460 , n31170 , n6249 );
    and g3137 ( n2399 , n17502 , n24295 );
    not g3138 ( n22673 , n25837 );
    xnor g3139 ( n22852 , n18563 , n12901 );
    xnor g3140 ( n26964 , n8175 , n27530 );
    not g3141 ( n3225 , n3613 );
    not g3142 ( n13391 , n6487 );
    not g3143 ( n6384 , n2687 );
    not g3144 ( n27775 , n28831 );
    xor g3145 ( n15941 , n19245 , n12931 );
    xnor g3146 ( n32020 , n5547 , n7736 );
    xnor g3147 ( n22582 , n18667 , n26082 );
    xnor g3148 ( n30 , n18609 , n26558 );
    or g3149 ( n24551 , n23934 , n11497 );
    or g3150 ( n27725 , n10496 , n14990 );
    xor g3151 ( n15505 , n7181 , n15742 );
    xor g3152 ( n14385 , n30919 , n12024 );
    xnor g3153 ( n6433 , n18531 , n499 );
    buf g3154 ( n19101 , n19177 );
    not g3155 ( n1817 , n6603 );
    and g3156 ( n8322 , n13320 , n27220 );
    not g3157 ( n15303 , n19187 );
    xnor g3158 ( n19542 , n25615 , n30246 );
    nor g3159 ( n3812 , n23306 , n20086 );
    not g3160 ( n11797 , n19356 );
    xnor g3161 ( n9075 , n10490 , n20038 );
    xnor g3162 ( n15608 , n15314 , n21836 );
    nor g3163 ( n15649 , n31845 , n5238 );
    not g3164 ( n5960 , n12056 );
    not g3165 ( n24365 , n9338 );
    or g3166 ( n23260 , n16272 , n31753 );
    nor g3167 ( n3694 , n30383 , n7193 );
    not g3168 ( n18345 , n9213 );
    xnor g3169 ( n30435 , n23140 , n7007 );
    or g3170 ( n28668 , n5789 , n17166 );
    xnor g3171 ( n14576 , n28201 , n5387 );
    or g3172 ( n566 , n2658 , n22252 );
    xnor g3173 ( n18159 , n13500 , n9134 );
    xnor g3174 ( n16789 , n10057 , n21138 );
    xnor g3175 ( n22040 , n6570 , n16830 );
    not g3176 ( n18059 , n25820 );
    and g3177 ( n3892 , n10201 , n31657 );
    or g3178 ( n30206 , n27321 , n21337 );
    not g3179 ( n20579 , n26299 );
    not g3180 ( n2736 , n18253 );
    not g3181 ( n24226 , n21997 );
    xnor g3182 ( n23081 , n10139 , n31060 );
    not g3183 ( n27525 , n7009 );
    not g3184 ( n20492 , n27550 );
    or g3185 ( n7886 , n20411 , n29789 );
    and g3186 ( n17075 , n17938 , n13662 );
    not g3187 ( n8410 , n2720 );
    or g3188 ( n15874 , n19264 , n24253 );
    xnor g3189 ( n20466 , n28053 , n20082 );
    xnor g3190 ( n22500 , n8062 , n8251 );
    not g3191 ( n12477 , n9706 );
    xor g3192 ( n14268 , n15002 , n12627 );
    and g3193 ( n14561 , n29724 , n146 );
    nor g3194 ( n7568 , n14795 , n18558 );
    xor g3195 ( n8775 , n7281 , n10204 );
    xnor g3196 ( n22106 , n4334 , n28870 );
    not g3197 ( n3568 , n3372 );
    xor g3198 ( n7619 , n4039 , n19289 );
    not g3199 ( n1499 , n28305 );
    not g3200 ( n18147 , n10949 );
    or g3201 ( n2118 , n24601 , n20718 );
    xnor g3202 ( n27211 , n2080 , n467 );
    and g3203 ( n12102 , n19789 , n17442 );
    xnor g3204 ( n8466 , n7603 , n20276 );
    and g3205 ( n4589 , n1912 , n15136 );
    not g3206 ( n7664 , n21964 );
    or g3207 ( n28138 , n5568 , n9507 );
    or g3208 ( n28140 , n34 , n116 );
    not g3209 ( n26982 , n10483 );
    not g3210 ( n20729 , n16406 );
    not g3211 ( n29513 , n7545 );
    not g3212 ( n18531 , n15121 );
    not g3213 ( n18768 , n15289 );
    or g3214 ( n27168 , n3004 , n22501 );
    buf g3215 ( n5077 , n17902 );
    and g3216 ( n26325 , n24972 , n28394 );
    not g3217 ( n629 , n23124 );
    not g3218 ( n31404 , n18305 );
    nor g3219 ( n18845 , n20139 , n6542 );
    xnor g3220 ( n12265 , n23465 , n2970 );
    and g3221 ( n22669 , n28443 , n8174 );
    and g3222 ( n31621 , n23191 , n24259 );
    not g3223 ( n30198 , n13707 );
    not g3224 ( n18711 , n3795 );
    xnor g3225 ( n17269 , n20878 , n15558 );
    xnor g3226 ( n9034 , n31787 , n3363 );
    nor g3227 ( n10556 , n28081 , n20920 );
    not g3228 ( n3354 , n5067 );
    or g3229 ( n14350 , n15727 , n24719 );
    or g3230 ( n21426 , n8368 , n10603 );
    not g3231 ( n24015 , n567 );
    not g3232 ( n12987 , n13260 );
    or g3233 ( n7079 , n29648 , n9810 );
    and g3234 ( n11420 , n23142 , n12887 );
    or g3235 ( n23392 , n6648 , n11164 );
    xnor g3236 ( n20561 , n20087 , n11792 );
    xnor g3237 ( n29206 , n1809 , n31343 );
    not g3238 ( n22004 , n3971 );
    or g3239 ( n17905 , n1597 , n19899 );
    nor g3240 ( n26188 , n6372 , n6393 );
    nor g3241 ( n20469 , n22422 , n14390 );
    not g3242 ( n18781 , n20225 );
    and g3243 ( n11156 , n6157 , n2729 );
    xnor g3244 ( n2333 , n19845 , n6036 );
    not g3245 ( n25405 , n31350 );
    xnor g3246 ( n29289 , n12619 , n7728 );
    not g3247 ( n10042 , n1722 );
    xnor g3248 ( n10355 , n11476 , n24160 );
    xnor g3249 ( n6711 , n20153 , n18052 );
    or g3250 ( n30743 , n1722 , n30999 );
    not g3251 ( n2597 , n11472 );
    not g3252 ( n30281 , n27368 );
    not g3253 ( n852 , n4085 );
    not g3254 ( n28843 , n27199 );
    or g3255 ( n8140 , n6306 , n3427 );
    nor g3256 ( n29366 , n31262 , n27128 );
    xnor g3257 ( n21743 , n27425 , n24634 );
    and g3258 ( n23422 , n15256 , n22178 );
    nor g3259 ( n22808 , n1039 , n14523 );
    not g3260 ( n30932 , n13225 );
    and g3261 ( n13314 , n25217 , n9800 );
    not g3262 ( n3095 , n105 );
    xnor g3263 ( n7875 , n27272 , n5685 );
    not g3264 ( n13989 , n7087 );
    not g3265 ( n24425 , n23496 );
    xor g3266 ( n8670 , n8189 , n5251 );
    not g3267 ( n10516 , n9475 );
    xnor g3268 ( n31050 , n16186 , n4365 );
    or g3269 ( n31118 , n30467 , n24881 );
    nor g3270 ( n14220 , n26414 , n6666 );
    not g3271 ( n5017 , n5985 );
    not g3272 ( n18077 , n25531 );
    or g3273 ( n8405 , n29203 , n6421 );
    xnor g3274 ( n27092 , n26473 , n11482 );
    and g3275 ( n27771 , n10571 , n1958 );
    nor g3276 ( n2654 , n28894 , n17737 );
    or g3277 ( n3397 , n14108 , n14740 );
    or g3278 ( n25456 , n5444 , n28798 );
    xnor g3279 ( n19885 , n24577 , n21718 );
    or g3280 ( n16700 , n16422 , n8116 );
    xnor g3281 ( n22449 , n24430 , n11279 );
    not g3282 ( n19668 , n14634 );
    and g3283 ( n2708 , n14857 , n13261 );
    not g3284 ( n16350 , n31698 );
    xnor g3285 ( n26090 , n20873 , n5962 );
    xnor g3286 ( n13536 , n29130 , n30670 );
    and g3287 ( n16838 , n21081 , n13306 );
    or g3288 ( n8884 , n5066 , n17915 );
    or g3289 ( n6752 , n16984 , n24001 );
    xnor g3290 ( n18399 , n26541 , n6603 );
    xnor g3291 ( n31353 , n31296 , n22211 );
    nor g3292 ( n3078 , n26259 , n15288 );
    not g3293 ( n3932 , n22747 );
    not g3294 ( n24914 , n11394 );
    xnor g3295 ( n21765 , n14132 , n24525 );
    nor g3296 ( n26309 , n16533 , n24992 );
    xnor g3297 ( n16604 , n1438 , n27939 );
    and g3298 ( n6724 , n1645 , n29554 );
    not g3299 ( n17429 , n11123 );
    and g3300 ( n29731 , n6759 , n19798 );
    not g3301 ( n19348 , n26733 );
    and g3302 ( n7201 , n21541 , n18716 );
    and g3303 ( n14154 , n7 , n1314 );
    xnor g3304 ( n14434 , n3697 , n5739 );
    or g3305 ( n10995 , n7414 , n14290 );
    not g3306 ( n15435 , n19312 );
    not g3307 ( n26552 , n19062 );
    and g3308 ( n15131 , n25423 , n7468 );
    not g3309 ( n16560 , n24712 );
    or g3310 ( n23084 , n29569 , n22331 );
    not g3311 ( n24302 , n5193 );
    and g3312 ( n31412 , n9671 , n6382 );
    not g3313 ( n20647 , n27213 );
    or g3314 ( n31449 , n7224 , n24353 );
    not g3315 ( n15472 , n16793 );
    or g3316 ( n18505 , n1549 , n9366 );
    and g3317 ( n5097 , n31378 , n9558 );
    not g3318 ( n12722 , n8616 );
    not g3319 ( n2137 , n17428 );
    xnor g3320 ( n7086 , n195 , n26926 );
    xnor g3321 ( n4886 , n22859 , n28752 );
    and g3322 ( n12470 , n19139 , n28771 );
    xor g3323 ( n2686 , n1474 , n1727 );
    xnor g3324 ( n23330 , n3601 , n26849 );
    or g3325 ( n4307 , n4207 , n7419 );
    or g3326 ( n8036 , n28363 , n31803 );
    and g3327 ( n18301 , n14500 , n26861 );
    and g3328 ( n19696 , n2072 , n2308 );
    or g3329 ( n30839 , n9045 , n23920 );
    or g3330 ( n6075 , n1563 , n20949 );
    and g3331 ( n13862 , n28380 , n28732 );
    not g3332 ( n21566 , n12649 );
    xnor g3333 ( n720 , n26954 , n26674 );
    not g3334 ( n5105 , n18979 );
    or g3335 ( n1393 , n31517 , n22378 );
    or g3336 ( n5049 , n11771 , n18345 );
    xnor g3337 ( n8309 , n27126 , n31773 );
    buf g3338 ( n19743 , n21748 );
    not g3339 ( n29432 , n10769 );
    nor g3340 ( n7571 , n30411 , n16134 );
    or g3341 ( n18495 , n31773 , n17308 );
    or g3342 ( n31987 , n1366 , n6725 );
    xnor g3343 ( n16052 , n4964 , n29132 );
    or g3344 ( n21214 , n6147 , n23742 );
    and g3345 ( n18440 , n25919 , n6033 );
    xnor g3346 ( n18245 , n21952 , n30079 );
    not g3347 ( n9684 , n14995 );
    not g3348 ( n5487 , n18467 );
    or g3349 ( n25292 , n26665 , n10755 );
    and g3350 ( n11167 , n17972 , n19136 );
    not g3351 ( n17644 , n27409 );
    not g3352 ( n25801 , n23097 );
    xnor g3353 ( n24991 , n28592 , n29390 );
    not g3354 ( n20781 , n3656 );
    xnor g3355 ( n11927 , n27633 , n18882 );
    or g3356 ( n18306 , n12503 , n3368 );
    xnor g3357 ( n16229 , n4031 , n30685 );
    not g3358 ( n30020 , n11588 );
    or g3359 ( n24101 , n24137 , n10443 );
    and g3360 ( n5198 , n7195 , n9090 );
    not g3361 ( n24151 , n4446 );
    or g3362 ( n24835 , n1891 , n27151 );
    xnor g3363 ( n24633 , n30275 , n12221 );
    nor g3364 ( n17703 , n30555 , n4990 );
    or g3365 ( n27568 , n9619 , n5988 );
    not g3366 ( n31324 , n18873 );
    not g3367 ( n11718 , n12409 );
    or g3368 ( n20112 , n14751 , n18804 );
    and g3369 ( n13238 , n18720 , n28576 );
    not g3370 ( n14869 , n19575 );
    or g3371 ( n13740 , n18572 , n20035 );
    xnor g3372 ( n31334 , n9932 , n6630 );
    or g3373 ( n2367 , n20250 , n5928 );
    xnor g3374 ( n19651 , n9313 , n24850 );
    xnor g3375 ( n21682 , n30525 , n18518 );
    or g3376 ( n24516 , n4815 , n980 );
    not g3377 ( n8724 , n22717 );
    or g3378 ( n24462 , n19303 , n27234 );
    or g3379 ( n3627 , n6218 , n16335 );
    or g3380 ( n31443 , n18145 , n3826 );
    xnor g3381 ( n21772 , n20856 , n2453 );
    or g3382 ( n13053 , n22692 , n16014 );
    or g3383 ( n1271 , n17639 , n16717 );
    nor g3384 ( n29592 , n10198 , n9078 );
    or g3385 ( n648 , n28912 , n17754 );
    and g3386 ( n3673 , n16566 , n3575 );
    nor g3387 ( n9386 , n20837 , n18725 );
    and g3388 ( n23677 , n11562 , n18932 );
    not g3389 ( n4490 , n19891 );
    not g3390 ( n3235 , n6695 );
    not g3391 ( n20578 , n5180 );
    not g3392 ( n3654 , n14925 );
    and g3393 ( n22370 , n6640 , n27426 );
    xnor g3394 ( n25297 , n2825 , n19217 );
    or g3395 ( n7082 , n15866 , n8091 );
    xnor g3396 ( n28166 , n17165 , n28559 );
    xnor g3397 ( n4409 , n8661 , n16240 );
    not g3398 ( n12962 , n13232 );
    xnor g3399 ( n8856 , n8928 , n209 );
    not g3400 ( n17130 , n4054 );
    xnor g3401 ( n72 , n9180 , n25555 );
    not g3402 ( n12629 , n6494 );
    xnor g3403 ( n21906 , n9565 , n30688 );
    nor g3404 ( n20623 , n16391 , n3426 );
    or g3405 ( n26685 , n3978 , n23495 );
    xnor g3406 ( n23555 , n28357 , n8398 );
    or g3407 ( n6741 , n42 , n25366 );
    or g3408 ( n11877 , n22104 , n21227 );
    not g3409 ( n31853 , n16925 );
    xnor g3410 ( n20811 , n26867 , n3858 );
    xnor g3411 ( n1413 , n8759 , n10629 );
    not g3412 ( n29683 , n9961 );
    xnor g3413 ( n2970 , n6117 , n29951 );
    not g3414 ( n4605 , n3614 );
    or g3415 ( n5842 , n3354 , n7442 );
    and g3416 ( n15407 , n22098 , n13372 );
    or g3417 ( n24756 , n21570 , n19802 );
    nor g3418 ( n11575 , n16803 , n10393 );
    and g3419 ( n19335 , n14358 , n5185 );
    not g3420 ( n29871 , n16264 );
    nor g3421 ( n4664 , n8042 , n28440 );
    and g3422 ( n14505 , n14820 , n26077 );
    and g3423 ( n1394 , n17416 , n13993 );
    or g3424 ( n23688 , n13484 , n1795 );
    and g3425 ( n27893 , n18038 , n11771 );
    or g3426 ( n28969 , n3984 , n5695 );
    xnor g3427 ( n10095 , n7074 , n15848 );
    or g3428 ( n16464 , n25369 , n6696 );
    and g3429 ( n18158 , n3897 , n8099 );
    not g3430 ( n18194 , n29604 );
    or g3431 ( n21953 , n31963 , n17909 );
    or g3432 ( n5505 , n18203 , n26977 );
    or g3433 ( n7472 , n2825 , n27930 );
    xnor g3434 ( n27483 , n31245 , n21098 );
    or g3435 ( n2452 , n7145 , n25139 );
    nor g3436 ( n22298 , n29059 , n1993 );
    not g3437 ( n22882 , n10169 );
    xnor g3438 ( n17438 , n31585 , n23927 );
    not g3439 ( n1225 , n17059 );
    nor g3440 ( n29784 , n11373 , n21551 );
    not g3441 ( n18743 , n26669 );
    or g3442 ( n10292 , n24932 , n31145 );
    and g3443 ( n19201 , n29864 , n21746 );
    not g3444 ( n7108 , n28818 );
    nor g3445 ( n6142 , n5616 , n18559 );
    nor g3446 ( n21484 , n15038 , n28370 );
    not g3447 ( n20798 , n18257 );
    not g3448 ( n14899 , n5688 );
    xnor g3449 ( n18903 , n20076 , n16911 );
    xnor g3450 ( n20860 , n28159 , n13318 );
    not g3451 ( n542 , n25730 );
    nor g3452 ( n16548 , n8163 , n3362 );
    nor g3453 ( n17421 , n27667 , n5710 );
    not g3454 ( n27120 , n7854 );
    not g3455 ( n167 , n25196 );
    and g3456 ( n301 , n14407 , n29783 );
    or g3457 ( n13664 , n13954 , n14343 );
    not g3458 ( n6126 , n31438 );
    nor g3459 ( n15540 , n30874 , n13447 );
    or g3460 ( n18642 , n23548 , n26432 );
    or g3461 ( n25959 , n26174 , n28788 );
    or g3462 ( n10571 , n21805 , n18315 );
    xnor g3463 ( n2869 , n11743 , n30706 );
    and g3464 ( n19799 , n11597 , n19887 );
    or g3465 ( n923 , n10118 , n30380 );
    not g3466 ( n13754 , n26279 );
    not g3467 ( n31917 , n5387 );
    not g3468 ( n15425 , n23829 );
    and g3469 ( n23606 , n3555 , n11429 );
    nor g3470 ( n20523 , n18733 , n10246 );
    not g3471 ( n17405 , n16856 );
    and g3472 ( n1148 , n15510 , n11863 );
    and g3473 ( n27675 , n26936 , n15725 );
    or g3474 ( n2699 , n468 , n2379 );
    xnor g3475 ( n18988 , n8986 , n6888 );
    or g3476 ( n12702 , n8781 , n16147 );
    xnor g3477 ( n25359 , n18355 , n12385 );
    xnor g3478 ( n8214 , n26641 , n22643 );
    and g3479 ( n14554 , n4605 , n2925 );
    or g3480 ( n14758 , n31835 , n27523 );
    xnor g3481 ( n7683 , n23770 , n19092 );
    or g3482 ( n11115 , n17981 , n27784 );
    xnor g3483 ( n24773 , n1559 , n14290 );
    xnor g3484 ( n6919 , n21367 , n29792 );
    not g3485 ( n24191 , n30756 );
    xnor g3486 ( n14074 , n6091 , n11217 );
    xor g3487 ( n9374 , n30616 , n23040 );
    xnor g3488 ( n4515 , n30932 , n1569 );
    and g3489 ( n11779 , n5310 , n16885 );
    xnor g3490 ( n26561 , n16988 , n25726 );
    not g3491 ( n11070 , n30614 );
    or g3492 ( n4112 , n5434 , n10530 );
    not g3493 ( n35 , n26824 );
    not g3494 ( n18501 , n24507 );
    xnor g3495 ( n30269 , n28369 , n20541 );
    xnor g3496 ( n18030 , n12939 , n29308 );
    not g3497 ( n24537 , n17493 );
    xor g3498 ( n30031 , n29105 , n10494 );
    not g3499 ( n16186 , n17382 );
    or g3500 ( n12132 , n25745 , n22522 );
    or g3501 ( n21092 , n24048 , n18885 );
    and g3502 ( n13788 , n6531 , n24665 );
    or g3503 ( n21843 , n3000 , n16887 );
    and g3504 ( n1607 , n3832 , n29122 );
    not g3505 ( n31631 , n7219 );
    not g3506 ( n26713 , n12246 );
    and g3507 ( n7620 , n30104 , n13879 );
    xnor g3508 ( n29576 , n10312 , n1670 );
    or g3509 ( n3687 , n7507 , n12523 );
    and g3510 ( n22986 , n22488 , n12956 );
    or g3511 ( n18043 , n22823 , n29749 );
    nor g3512 ( n26777 , n3366 , n11773 );
    not g3513 ( n16637 , n24901 );
    nor g3514 ( n5289 , n27444 , n16492 );
    not g3515 ( n8936 , n21326 );
    and g3516 ( n30044 , n24742 , n5010 );
    and g3517 ( n10100 , n27450 , n28733 );
    and g3518 ( n16640 , n14546 , n18901 );
    or g3519 ( n21709 , n23294 , n4022 );
    not g3520 ( n26174 , n5147 );
    not g3521 ( n15772 , n18487 );
    not g3522 ( n3548 , n31324 );
    nor g3523 ( n11278 , n30245 , n13797 );
    not g3524 ( n14458 , n2588 );
    and g3525 ( n11710 , n12331 , n18194 );
    not g3526 ( n31963 , n11738 );
    xnor g3527 ( n6396 , n12473 , n2357 );
    or g3528 ( n10644 , n26296 , n10272 );
    not g3529 ( n23562 , n10532 );
    nor g3530 ( n22240 , n29095 , n4489 );
    xnor g3531 ( n11811 , n23484 , n29967 );
    not g3532 ( n30018 , n2122 );
    not g3533 ( n18275 , n16982 );
    nor g3534 ( n4811 , n1819 , n7218 );
    not g3535 ( n3581 , n19127 );
    xnor g3536 ( n23706 , n27885 , n26996 );
    nor g3537 ( n11988 , n27850 , n1919 );
    xor g3538 ( n12175 , n9699 , n13700 );
    nor g3539 ( n5538 , n16587 , n31182 );
    and g3540 ( n4058 , n3960 , n11265 );
    not g3541 ( n9039 , n6511 );
    xnor g3542 ( n4368 , n24192 , n19274 );
    not g3543 ( n17516 , n13864 );
    and g3544 ( n29755 , n6220 , n2304 );
    xnor g3545 ( n27342 , n204 , n22712 );
    not g3546 ( n10301 , n16778 );
    or g3547 ( n14023 , n12959 , n30813 );
    and g3548 ( n8835 , n4966 , n22136 );
    nor g3549 ( n26018 , n15873 , n4939 );
    not g3550 ( n6926 , n25994 );
    or g3551 ( n26334 , n10286 , n8231 );
    xor g3552 ( n15798 , n6051 , n8240 );
    or g3553 ( n7437 , n28828 , n11852 );
    xnor g3554 ( n30025 , n6262 , n8213 );
    not g3555 ( n10104 , n775 );
    or g3556 ( n28125 , n12998 , n5876 );
    not g3557 ( n1113 , n28205 );
    not g3558 ( n16452 , n22170 );
    not g3559 ( n3262 , n4297 );
    not g3560 ( n5417 , n17515 );
    not g3561 ( n16368 , n14630 );
    xnor g3562 ( n25053 , n19279 , n14567 );
    not g3563 ( n16319 , n12082 );
    not g3564 ( n1072 , n9512 );
    nor g3565 ( n3102 , n9146 , n335 );
    or g3566 ( n2471 , n19366 , n13041 );
    not g3567 ( n13972 , n19255 );
    nor g3568 ( n12504 , n27974 , n10185 );
    not g3569 ( n1488 , n7876 );
    nor g3570 ( n25692 , n25527 , n17302 );
    nor g3571 ( n31648 , n9788 , n4714 );
    and g3572 ( n11408 , n24882 , n21145 );
    or g3573 ( n24802 , n6553 , n30035 );
    xnor g3574 ( n26237 , n19826 , n5416 );
    xnor g3575 ( n7634 , n31910 , n16308 );
    not g3576 ( n12694 , n17851 );
    or g3577 ( n9671 , n18142 , n18436 );
    xnor g3578 ( n14137 , n29942 , n3352 );
    or g3579 ( n22404 , n31452 , n15626 );
    not g3580 ( n21325 , n30182 );
    not g3581 ( n9579 , n25042 );
    not g3582 ( n25950 , n5022 );
    xnor g3583 ( n7847 , n22759 , n22868 );
    not g3584 ( n16625 , n15382 );
    nor g3585 ( n5955 , n31591 , n26525 );
    or g3586 ( n11732 , n138 , n19042 );
    or g3587 ( n19766 , n26084 , n22080 );
    or g3588 ( n9732 , n4895 , n214 );
    not g3589 ( n826 , n13507 );
    xnor g3590 ( n19998 , n20495 , n6331 );
    not g3591 ( n315 , n2509 );
    xnor g3592 ( n6592 , n13083 , n823 );
    not g3593 ( n16982 , n2185 );
    not g3594 ( n18969 , n2727 );
    not g3595 ( n2329 , n10911 );
    nor g3596 ( n25071 , n27183 , n14586 );
    or g3597 ( n28079 , n16560 , n21033 );
    nor g3598 ( n22338 , n16195 , n24483 );
    xnor g3599 ( n1123 , n30096 , n25889 );
    nor g3600 ( n20024 , n23834 , n9826 );
    xor g3601 ( n22935 , n22214 , n2615 );
    nor g3602 ( n1408 , n31313 , n20153 );
    not g3603 ( n1537 , n31688 );
    xnor g3604 ( n28458 , n31756 , n15820 );
    and g3605 ( n844 , n21837 , n18539 );
    or g3606 ( n28889 , n24421 , n774 );
    nor g3607 ( n12708 , n1692 , n33 );
    not g3608 ( n22748 , n8600 );
    not g3609 ( n14423 , n31095 );
    not g3610 ( n28574 , n24306 );
    or g3611 ( n16432 , n23700 , n27036 );
    not g3612 ( n4434 , n1879 );
    not g3613 ( n28633 , n18555 );
    or g3614 ( n27526 , n28080 , n22583 );
    xnor g3615 ( n21266 , n13496 , n17635 );
    or g3616 ( n15021 , n21310 , n15613 );
    and g3617 ( n26048 , n21190 , n20566 );
    or g3618 ( n31089 , n24521 , n151 );
    xnor g3619 ( n2290 , n12894 , n13164 );
    xnor g3620 ( n9551 , n25523 , n15945 );
    or g3621 ( n17529 , n3178 , n23446 );
    and g3622 ( n10295 , n3395 , n13846 );
    nor g3623 ( n31681 , n19058 , n6496 );
    nor g3624 ( n25870 , n27533 , n6030 );
    and g3625 ( n18160 , n4880 , n3414 );
    nor g3626 ( n24412 , n14186 , n11642 );
    nor g3627 ( n21062 , n11610 , n31252 );
    xnor g3628 ( n25790 , n31201 , n20880 );
    not g3629 ( n16457 , n10082 );
    nor g3630 ( n16630 , n10729 , n14214 );
    xnor g3631 ( n3976 , n25798 , n30593 );
    not g3632 ( n19695 , n1203 );
    nor g3633 ( n20524 , n26974 , n16986 );
    not g3634 ( n15204 , n7184 );
    and g3635 ( n1634 , n17407 , n26783 );
    and g3636 ( n5354 , n31994 , n10446 );
    not g3637 ( n22497 , n14388 );
    and g3638 ( n5383 , n28715 , n13711 );
    or g3639 ( n18497 , n7506 , n19335 );
    not g3640 ( n5250 , n30951 );
    not g3641 ( n275 , n17803 );
    and g3642 ( n24170 , n21283 , n12977 );
    nor g3643 ( n27224 , n14330 , n16416 );
    xnor g3644 ( n29456 , n22817 , n31199 );
    not g3645 ( n4511 , n2001 );
    xnor g3646 ( n931 , n28356 , n12143 );
    or g3647 ( n18822 , n3552 , n17078 );
    or g3648 ( n13340 , n18681 , n24965 );
    xnor g3649 ( n5329 , n17016 , n6196 );
    or g3650 ( n22391 , n28450 , n16366 );
    not g3651 ( n11007 , n5300 );
    or g3652 ( n2611 , n10712 , n14145 );
    xnor g3653 ( n7511 , n6685 , n20452 );
    or g3654 ( n1060 , n14369 , n5830 );
    not g3655 ( n18067 , n31326 );
    and g3656 ( n26295 , n30524 , n20309 );
    and g3657 ( n26274 , n29612 , n4139 );
    nor g3658 ( n2697 , n27829 , n14503 );
    and g3659 ( n13443 , n155 , n12565 );
    nor g3660 ( n20470 , n10106 , n31860 );
    xnor g3661 ( n5531 , n20003 , n29057 );
    or g3662 ( n31273 , n9954 , n27628 );
    or g3663 ( n17412 , n11347 , n30154 );
    not g3664 ( n15683 , n21192 );
    not g3665 ( n10614 , n26269 );
    or g3666 ( n19638 , n18018 , n13426 );
    or g3667 ( n24720 , n5044 , n6134 );
    not g3668 ( n1351 , n18850 );
    not g3669 ( n16182 , n23400 );
    and g3670 ( n1919 , n19767 , n12531 );
    xnor g3671 ( n20185 , n11132 , n17995 );
    or g3672 ( n9020 , n23027 , n11917 );
    xnor g3673 ( n10511 , n29420 , n30982 );
    and g3674 ( n26637 , n8957 , n6225 );
    not g3675 ( n10223 , n7623 );
    not g3676 ( n21785 , n28044 );
    xnor g3677 ( n1924 , n10521 , n25089 );
    xnor g3678 ( n3466 , n12072 , n17019 );
    xnor g3679 ( n20274 , n25111 , n25500 );
    xnor g3680 ( n7231 , n26357 , n8696 );
    xnor g3681 ( n31515 , n28768 , n31309 );
    and g3682 ( n21333 , n29497 , n23764 );
    and g3683 ( n9507 , n9440 , n15831 );
    xnor g3684 ( n30672 , n25016 , n16540 );
    and g3685 ( n4039 , n29925 , n11871 );
    and g3686 ( n2312 , n15749 , n24184 );
    not g3687 ( n1711 , n4221 );
    not g3688 ( n29567 , n8622 );
    xnor g3689 ( n13814 , n15412 , n11845 );
    or g3690 ( n1644 , n13855 , n15669 );
    xor g3691 ( n21954 , n17860 , n8435 );
    and g3692 ( n16595 , n21274 , n12253 );
    buf g3693 ( n8901 , n31356 );
    and g3694 ( n17414 , n2625 , n18207 );
    nor g3695 ( n17856 , n23843 , n21007 );
    or g3696 ( n9991 , n8975 , n30536 );
    and g3697 ( n23629 , n26702 , n27600 );
    not g3698 ( n9743 , n13451 );
    xnor g3699 ( n5896 , n24343 , n3281 );
    not g3700 ( n23490 , n5165 );
    and g3701 ( n18263 , n13611 , n2860 );
    xnor g3702 ( n20960 , n11382 , n5680 );
    not g3703 ( n9543 , n19336 );
    nor g3704 ( n16758 , n1529 , n20667 );
    not g3705 ( n10870 , n21007 );
    nor g3706 ( n15016 , n17585 , n20486 );
    xnor g3707 ( n18293 , n15664 , n8718 );
    nor g3708 ( n960 , n24095 , n17831 );
    xnor g3709 ( n10951 , n19598 , n28207 );
    nor g3710 ( n8523 , n8714 , n13908 );
    or g3711 ( n2940 , n9414 , n28022 );
    not g3712 ( n19240 , n2677 );
    or g3713 ( n1092 , n9255 , n1133 );
    not g3714 ( n11513 , n19625 );
    xnor g3715 ( n4095 , n29585 , n23409 );
    or g3716 ( n11311 , n27291 , n7416 );
    nor g3717 ( n19374 , n14777 , n17670 );
    and g3718 ( n14395 , n16503 , n15508 );
    or g3719 ( n8883 , n11989 , n16479 );
    xnor g3720 ( n9675 , n30301 , n15714 );
    and g3721 ( n1544 , n24825 , n991 );
    and g3722 ( n19664 , n18546 , n2598 );
    or g3723 ( n13965 , n29471 , n17826 );
    and g3724 ( n29482 , n24868 , n18879 );
    xnor g3725 ( n7095 , n4992 , n31722 );
    xnor g3726 ( n10860 , n5731 , n19663 );
    or g3727 ( n11633 , n5365 , n20809 );
    xnor g3728 ( n7882 , n22673 , n22077 );
    nor g3729 ( n1505 , n11577 , n6230 );
    xnor g3730 ( n17920 , n9469 , n29569 );
    and g3731 ( n2551 , n698 , n22886 );
    xnor g3732 ( n18473 , n9528 , n12609 );
    xnor g3733 ( n1428 , n4738 , n26999 );
    or g3734 ( n4101 , n23121 , n21751 );
    nor g3735 ( n6476 , n30405 , n18403 );
    and g3736 ( n31588 , n15919 , n19203 );
    xnor g3737 ( n17607 , n407 , n92 );
    or g3738 ( n14138 , n14213 , n27288 );
    xnor g3739 ( n29316 , n11588 , n5326 );
    and g3740 ( n20132 , n20736 , n30936 );
    not g3741 ( n1172 , n26830 );
    and g3742 ( n18426 , n28167 , n15728 );
    or g3743 ( n5283 , n19132 , n16598 );
    not g3744 ( n7140 , n13663 );
    not g3745 ( n4226 , n29721 );
    not g3746 ( n22428 , n22882 );
    or g3747 ( n15564 , n30047 , n22552 );
    or g3748 ( n10215 , n31276 , n322 );
    xnor g3749 ( n27226 , n13945 , n27344 );
    xnor g3750 ( n25524 , n2344 , n3630 );
    and g3751 ( n24467 , n18551 , n21136 );
    and g3752 ( n21620 , n71 , n11661 );
    and g3753 ( n7848 , n25958 , n5948 );
    and g3754 ( n1688 , n17040 , n26339 );
    not g3755 ( n22543 , n15041 );
    xnor g3756 ( n32007 , n3402 , n19397 );
    xnor g3757 ( n26834 , n5514 , n5420 );
    or g3758 ( n29258 , n3553 , n5586 );
    not g3759 ( n31731 , n9228 );
    not g3760 ( n7560 , n22429 );
    and g3761 ( n31684 , n17311 , n6444 );
    not g3762 ( n16678 , n3495 );
    and g3763 ( n7020 , n5084 , n3044 );
    nor g3764 ( n7913 , n1000 , n18486 );
    xnor g3765 ( n11428 , n2568 , n6615 );
    or g3766 ( n16846 , n5500 , n2439 );
    or g3767 ( n9013 , n11462 , n9461 );
    not g3768 ( n9901 , n31102 );
    xnor g3769 ( n12944 , n1426 , n14975 );
    xnor g3770 ( n1982 , n27355 , n19274 );
    xnor g3771 ( n4987 , n28385 , n28643 );
    and g3772 ( n12033 , n22805 , n5196 );
    nor g3773 ( n14981 , n28183 , n14438 );
    not g3774 ( n20174 , n8110 );
    xnor g3775 ( n15147 , n2145 , n16411 );
    not g3776 ( n24324 , n10310 );
    nor g3777 ( n5218 , n7261 , n16282 );
    or g3778 ( n17433 , n16015 , n12415 );
    not g3779 ( n4737 , n17219 );
    or g3780 ( n29627 , n26344 , n7326 );
    nor g3781 ( n5583 , n30002 , n29471 );
    or g3782 ( n4485 , n8988 , n26373 );
    xnor g3783 ( n16120 , n7887 , n8455 );
    or g3784 ( n1303 , n12536 , n14210 );
    not g3785 ( n29766 , n28767 );
    nor g3786 ( n28100 , n12221 , n30433 );
    xnor g3787 ( n10254 , n23781 , n1255 );
    and g3788 ( n22417 , n21479 , n15537 );
    or g3789 ( n6004 , n8025 , n18526 );
    or g3790 ( n16831 , n9468 , n7123 );
    xnor g3791 ( n30904 , n8060 , n28918 );
    xnor g3792 ( n16953 , n12225 , n30367 );
    xnor g3793 ( n19055 , n4910 , n3485 );
    and g3794 ( n9657 , n16280 , n23956 );
    nor g3795 ( n5213 , n6071 , n6740 );
    xnor g3796 ( n30005 , n27681 , n20002 );
    or g3797 ( n4705 , n29142 , n30263 );
    xnor g3798 ( n6988 , n26773 , n20203 );
    not g3799 ( n21506 , n21369 );
    xnor g3800 ( n9853 , n24566 , n252 );
    or g3801 ( n17528 , n12430 , n28923 );
    or g3802 ( n1706 , n6657 , n16777 );
    xnor g3803 ( n20931 , n23860 , n3419 );
    not g3804 ( n15620 , n26004 );
    or g3805 ( n6572 , n14341 , n19112 );
    not g3806 ( n30195 , n6180 );
    xnor g3807 ( n5944 , n29140 , n11584 );
    not g3808 ( n11248 , n780 );
    xnor g3809 ( n13289 , n19075 , n22182 );
    not g3810 ( n21495 , n10790 );
    nor g3811 ( n6837 , n10433 , n23547 );
    and g3812 ( n16739 , n17488 , n8450 );
    xor g3813 ( n6100 , n25385 , n23521 );
    xnor g3814 ( n31965 , n9004 , n27517 );
    xor g3815 ( n10904 , n30082 , n306 );
    not g3816 ( n15714 , n10129 );
    or g3817 ( n10882 , n16782 , n5159 );
    or g3818 ( n18717 , n15622 , n29893 );
    not g3819 ( n10863 , n9835 );
    or g3820 ( n11091 , n21104 , n23932 );
    not g3821 ( n28437 , n23868 );
    or g3822 ( n2418 , n7374 , n26922 );
    not g3823 ( n11052 , n18512 );
    or g3824 ( n4346 , n17149 , n3131 );
    xnor g3825 ( n6356 , n17632 , n31419 );
    not g3826 ( n9690 , n856 );
    not g3827 ( n15975 , n27805 );
    xnor g3828 ( n25716 , n24025 , n20591 );
    not g3829 ( n22754 , n12779 );
    and g3830 ( n7102 , n7432 , n28156 );
    not g3831 ( n1913 , n20453 );
    or g3832 ( n19411 , n4557 , n24505 );
    and g3833 ( n25168 , n31747 , n19602 );
    and g3834 ( n30750 , n18864 , n4580 );
    or g3835 ( n3925 , n17337 , n26314 );
    nor g3836 ( n26280 , n27008 , n4050 );
    not g3837 ( n26024 , n12498 );
    nor g3838 ( n31974 , n24991 , n18691 );
    and g3839 ( n10540 , n20901 , n27626 );
    or g3840 ( n3779 , n25917 , n29614 );
    not g3841 ( n16514 , n8720 );
    or g3842 ( n6922 , n28326 , n27764 );
    or g3843 ( n17594 , n11262 , n31248 );
    and g3844 ( n7792 , n18196 , n13056 );
    and g3845 ( n19526 , n19844 , n31436 );
    not g3846 ( n206 , n13059 );
    not g3847 ( n28356 , n10114 );
    xnor g3848 ( n27510 , n6997 , n16393 );
    and g3849 ( n610 , n15186 , n9941 );
    and g3850 ( n5700 , n10590 , n12578 );
    not g3851 ( n19299 , n17257 );
    or g3852 ( n15905 , n8474 , n22489 );
    not g3853 ( n158 , n8526 );
    and g3854 ( n5129 , n2474 , n28660 );
    xnor g3855 ( n31317 , n31816 , n8028 );
    not g3856 ( n27889 , n27579 );
    or g3857 ( n11530 , n4429 , n31075 );
    xnor g3858 ( n6602 , n31997 , n12577 );
    or g3859 ( n18770 , n6516 , n31768 );
    not g3860 ( n15387 , n27153 );
    xnor g3861 ( n15045 , n2865 , n5817 );
    not g3862 ( n29025 , n23438 );
    or g3863 ( n17408 , n26252 , n1909 );
    xnor g3864 ( n31545 , n5940 , n28113 );
    and g3865 ( n7303 , n12044 , n11780 );
    not g3866 ( n5319 , n26213 );
    xnor g3867 ( n29207 , n19414 , n31336 );
    not g3868 ( n24441 , n15213 );
    not g3869 ( n17004 , n22525 );
    xnor g3870 ( n26780 , n6152 , n24129 );
    or g3871 ( n26631 , n15181 , n30687 );
    or g3872 ( n27347 , n13183 , n5427 );
    not g3873 ( n28400 , n2973 );
    not g3874 ( n11680 , n13197 );
    not g3875 ( n12001 , n13635 );
    not g3876 ( n2086 , n12209 );
    nor g3877 ( n4927 , n14037 , n10939 );
    or g3878 ( n6894 , n10941 , n16899 );
    and g3879 ( n25926 , n758 , n2934 );
    not g3880 ( n2791 , n10508 );
    not g3881 ( n16057 , n31603 );
    and g3882 ( n26742 , n21236 , n9175 );
    xnor g3883 ( n27979 , n27801 , n10284 );
    not g3884 ( n5147 , n21633 );
    xnor g3885 ( n25734 , n138 , n10114 );
    xnor g3886 ( n27304 , n5741 , n27310 );
    not g3887 ( n2029 , n19837 );
    not g3888 ( n28790 , n2889 );
    and g3889 ( n20100 , n25898 , n27027 );
    xnor g3890 ( n17672 , n31523 , n10902 );
    not g3891 ( n16352 , n3545 );
    and g3892 ( n29464 , n11237 , n21690 );
    xnor g3893 ( n20098 , n25504 , n16302 );
    or g3894 ( n21541 , n22208 , n28868 );
    xnor g3895 ( n18128 , n29541 , n21994 );
    not g3896 ( n9387 , n31898 );
    not g3897 ( n21891 , n18251 );
    and g3898 ( n27145 , n27715 , n21136 );
    nor g3899 ( n5857 , n18655 , n26398 );
    not g3900 ( n23810 , n16155 );
    xnor g3901 ( n7921 , n4195 , n18449 );
    xnor g3902 ( n23758 , n27581 , n26541 );
    not g3903 ( n25931 , n5798 );
    not g3904 ( n10008 , n26179 );
    or g3905 ( n23267 , n2429 , n1052 );
    and g3906 ( n23548 , n21468 , n11672 );
    xnor g3907 ( n26388 , n7806 , n21502 );
    not g3908 ( n17072 , n23335 );
    xnor g3909 ( n30649 , n3666 , n8676 );
    or g3910 ( n20191 , n27478 , n30759 );
    xnor g3911 ( n29830 , n8178 , n17068 );
    or g3912 ( n20903 , n27612 , n17564 );
    not g3913 ( n255 , n23312 );
    nor g3914 ( n25567 , n13398 , n2717 );
    xnor g3915 ( n6778 , n22069 , n17959 );
    not g3916 ( n8328 , n1800 );
    xor g3917 ( n26809 , n15066 , n1234 );
    xnor g3918 ( n6082 , n28971 , n30164 );
    nor g3919 ( n9927 , n27453 , n12696 );
    xnor g3920 ( n24100 , n23682 , n24554 );
    and g3921 ( n4668 , n16540 , n28500 );
    xnor g3922 ( n12310 , n12299 , n21301 );
    and g3923 ( n30875 , n23001 , n17778 );
    not g3924 ( n19756 , n3359 );
    and g3925 ( n25533 , n19457 , n6719 );
    not g3926 ( n7957 , n29569 );
    not g3927 ( n13233 , n2693 );
    not g3928 ( n21720 , n26114 );
    not g3929 ( n21883 , n5881 );
    not g3930 ( n3454 , n11984 );
    xnor g3931 ( n23943 , n15333 , n24797 );
    xnor g3932 ( n1284 , n2282 , n763 );
    and g3933 ( n9315 , n16507 , n26099 );
    not g3934 ( n27270 , n30180 );
    and g3935 ( n16472 , n27812 , n30107 );
    or g3936 ( n307 , n1129 , n21338 );
    or g3937 ( n18163 , n11218 , n12349 );
    not g3938 ( n17379 , n16023 );
    and g3939 ( n5722 , n11040 , n19390 );
    xnor g3940 ( n11074 , n30276 , n15113 );
    not g3941 ( n22173 , n15674 );
    nor g3942 ( n6376 , n4130 , n19343 );
    xnor g3943 ( n3261 , n8903 , n5778 );
    nor g3944 ( n13575 , n508 , n31914 );
    nor g3945 ( n10041 , n2250 , n30812 );
    xnor g3946 ( n16795 , n12430 , n28695 );
    and g3947 ( n29602 , n16224 , n4064 );
    not g3948 ( n12992 , n24578 );
    not g3949 ( n17335 , n20857 );
    not g3950 ( n7433 , n5102 );
    xnor g3951 ( n13291 , n12444 , n24181 );
    or g3952 ( n26046 , n26734 , n26180 );
    and g3953 ( n6502 , n8265 , n28808 );
    and g3954 ( n19519 , n24310 , n26981 );
    not g3955 ( n18966 , n16651 );
    not g3956 ( n14119 , n757 );
    xnor g3957 ( n15020 , n11718 , n10114 );
    not g3958 ( n8283 , n2934 );
    not g3959 ( n30021 , n28028 );
    not g3960 ( n12502 , n10638 );
    xnor g3961 ( n7299 , n7022 , n5715 );
    nor g3962 ( n28802 , n18647 , n17941 );
    not g3963 ( n29669 , n27848 );
    not g3964 ( n12473 , n26436 );
    not g3965 ( n22587 , n28336 );
    or g3966 ( n30631 , n953 , n18530 );
    not g3967 ( n16859 , n3914 );
    or g3968 ( n455 , n31280 , n8926 );
    xnor g3969 ( n25781 , n17711 , n22531 );
    or g3970 ( n26572 , n31862 , n4876 );
    xnor g3971 ( n18544 , n13275 , n30651 );
    and g3972 ( n30767 , n22054 , n12393 );
    or g3973 ( n27119 , n26896 , n29860 );
    xnor g3974 ( n836 , n8350 , n15124 );
    not g3975 ( n31483 , n14477 );
    xor g3976 ( n26271 , n10755 , n12099 );
    xnor g3977 ( n14917 , n10643 , n26665 );
    not g3978 ( n4812 , n1616 );
    xnor g3979 ( n30414 , n18546 , n31740 );
    xnor g3980 ( n15520 , n4944 , n7217 );
    xnor g3981 ( n31079 , n18360 , n22665 );
    not g3982 ( n17862 , n15299 );
    xor g3983 ( n29445 , n29120 , n24221 );
    not g3984 ( n28906 , n5733 );
    xor g3985 ( n19185 , n15208 , n21301 );
    or g3986 ( n2478 , n3480 , n12639 );
    xnor g3987 ( n24127 , n2100 , n11028 );
    not g3988 ( n18318 , n13491 );
    not g3989 ( n15029 , n19013 );
    and g3990 ( n15788 , n15256 , n18559 );
    xnor g3991 ( n18887 , n9489 , n4630 );
    or g3992 ( n9356 , n10028 , n17482 );
    and g3993 ( n1182 , n18396 , n1449 );
    and g3994 ( n1313 , n9394 , n26135 );
    xnor g3995 ( n11433 , n1560 , n25359 );
    and g3996 ( n30915 , n17554 , n21120 );
    xor g3997 ( n23312 , n23117 , n31890 );
    xnor g3998 ( n15132 , n25867 , n11041 );
    and g3999 ( n10671 , n11973 , n14624 );
    not g4000 ( n3311 , n15027 );
    or g4001 ( n19634 , n1314 , n7194 );
    and g4002 ( n15567 , n16083 , n21956 );
    not g4003 ( n21439 , n19478 );
    nor g4004 ( n28388 , n12207 , n23184 );
    not g4005 ( n22738 , n8316 );
    xnor g4006 ( n3527 , n18391 , n3782 );
    or g4007 ( n18721 , n7897 , n21820 );
    and g4008 ( n21196 , n27673 , n8909 );
    or g4009 ( n15163 , n8956 , n959 );
    or g4010 ( n28086 , n17585 , n18312 );
    and g4011 ( n14 , n14376 , n24246 );
    or g4012 ( n15581 , n21381 , n19444 );
    xnor g4013 ( n17471 , n7429 , n14806 );
    and g4014 ( n13646 , n20815 , n22665 );
    nor g4015 ( n1026 , n14025 , n17024 );
    xnor g4016 ( n2129 , n15052 , n29888 );
    not g4017 ( n19340 , n26943 );
    nor g4018 ( n30312 , n19317 , n19652 );
    xnor g4019 ( n29454 , n15029 , n10322 );
    xnor g4020 ( n16077 , n1446 , n26400 );
    or g4021 ( n8624 , n30287 , n26749 );
    or g4022 ( n6744 , n9952 , n22767 );
    not g4023 ( n21337 , n513 );
    not g4024 ( n4255 , n13210 );
    xnor g4025 ( n28679 , n7566 , n3281 );
    not g4026 ( n31201 , n25202 );
    xnor g4027 ( n28852 , n15720 , n31869 );
    not g4028 ( n25880 , n25499 );
    nor g4029 ( n27203 , n29805 , n10486 );
    or g4030 ( n4840 , n15884 , n30988 );
    nor g4031 ( n4038 , n12125 , n27899 );
    xnor g4032 ( n18423 , n17373 , n22036 );
    or g4033 ( n27622 , n445 , n26114 );
    and g4034 ( n24307 , n23006 , n26883 );
    nor g4035 ( n14439 , n10239 , n4672 );
    nor g4036 ( n7889 , n6717 , n30218 );
    xnor g4037 ( n15826 , n16335 , n9797 );
    xnor g4038 ( n29650 , n8799 , n14582 );
    not g4039 ( n11130 , n22111 );
    and g4040 ( n28871 , n2222 , n26854 );
    xnor g4041 ( n14167 , n4351 , n14454 );
    and g4042 ( n14922 , n1352 , n19301 );
    or g4043 ( n16499 , n20573 , n8360 );
    and g4044 ( n17486 , n10520 , n11926 );
    and g4045 ( n19550 , n9967 , n12770 );
    not g4046 ( n18990 , n28417 );
    and g4047 ( n13810 , n20053 , n23351 );
    not g4048 ( n17730 , n30148 );
    not g4049 ( n2485 , n9580 );
    or g4050 ( n27063 , n18063 , n6198 );
    not g4051 ( n20538 , n10451 );
    xnor g4052 ( n7745 , n7890 , n8030 );
    and g4053 ( n26164 , n25663 , n3243 );
    not g4054 ( n25629 , n8201 );
    xnor g4055 ( n30757 , n23957 , n23142 );
    nor g4056 ( n28684 , n16151 , n18977 );
    nor g4057 ( n23116 , n10158 , n41 );
    xnor g4058 ( n22743 , n31220 , n24245 );
    xnor g4059 ( n8094 , n3904 , n12226 );
    not g4060 ( n4404 , n27452 );
    and g4061 ( n11893 , n11118 , n3050 );
    or g4062 ( n11715 , n14974 , n6754 );
    or g4063 ( n4800 , n11636 , n9788 );
    xnor g4064 ( n21774 , n19682 , n12435 );
    not g4065 ( n29600 , n1188 );
    nor g4066 ( n31675 , n9528 , n27916 );
    or g4067 ( n30876 , n1850 , n6057 );
    not g4068 ( n2800 , n28712 );
    not g4069 ( n643 , n14595 );
    xnor g4070 ( n20627 , n8035 , n10912 );
    or g4071 ( n31660 , n508 , n18764 );
    xnor g4072 ( n21250 , n2447 , n6141 );
    and g4073 ( n2496 , n26119 , n1117 );
    and g4074 ( n22462 , n27188 , n10783 );
    nor g4075 ( n30484 , n9480 , n15343 );
    xnor g4076 ( n27106 , n12950 , n29049 );
    not g4077 ( n11924 , n26725 );
    or g4078 ( n30563 , n11998 , n18710 );
    or g4079 ( n15747 , n21761 , n20757 );
    xnor g4080 ( n3224 , n18646 , n6961 );
    xnor g4081 ( n9113 , n28819 , n28615 );
    or g4082 ( n8823 , n15179 , n966 );
    xnor g4083 ( n14098 , n17488 , n27179 );
    xor g4084 ( n11445 , n13552 , n5388 );
    xnor g4085 ( n25043 , n19667 , n31802 );
    xor g4086 ( n5579 , n13142 , n24422 );
    xnor g4087 ( n26836 , n5314 , n23723 );
    nor g4088 ( n25654 , n31783 , n21494 );
    not g4089 ( n16381 , n19224 );
    or g4090 ( n7322 , n27218 , n7932 );
    not g4091 ( n17355 , n3486 );
    not g4092 ( n15457 , n10143 );
    or g4093 ( n12499 , n11931 , n14332 );
    and g4094 ( n28518 , n26468 , n18719 );
    nor g4095 ( n17716 , n22467 , n16038 );
    xnor g4096 ( n11521 , n19668 , n24322 );
    xnor g4097 ( n25192 , n26651 , n27150 );
    and g4098 ( n20280 , n26478 , n10245 );
    or g4099 ( n21203 , n4195 , n27117 );
    xnor g4100 ( n264 , n9469 , n22922 );
    not g4101 ( n6069 , n23455 );
    not g4102 ( n30392 , n1327 );
    or g4103 ( n25400 , n11256 , n22544 );
    not g4104 ( n967 , n3256 );
    xnor g4105 ( n2354 , n28480 , n5782 );
    xnor g4106 ( n214 , n11495 , n23138 );
    not g4107 ( n21556 , n12867 );
    nor g4108 ( n17956 , n29695 , n21491 );
    or g4109 ( n1469 , n19156 , n119 );
    xor g4110 ( n6938 , n19422 , n1616 );
    not g4111 ( n4796 , n21851 );
    xnor g4112 ( n16737 , n28312 , n20722 );
    not g4113 ( n17517 , n13397 );
    or g4114 ( n15395 , n12012 , n20349 );
    not g4115 ( n25512 , n28333 );
    xnor g4116 ( n23469 , n6318 , n15665 );
    or g4117 ( n31398 , n30612 , n1580 );
    or g4118 ( n9363 , n4104 , n17198 );
    and g4119 ( n30055 , n1364 , n20719 );
    or g4120 ( n25925 , n25078 , n12022 );
    and g4121 ( n8750 , n28143 , n16653 );
    or g4122 ( n28944 , n13224 , n11911 );
    not g4123 ( n14351 , n26308 );
    and g4124 ( n28062 , n18847 , n19990 );
    not g4125 ( n4334 , n1670 );
    nor g4126 ( n27610 , n11643 , n177 );
    and g4127 ( n1914 , n31298 , n15229 );
    and g4128 ( n22914 , n12043 , n14520 );
    not g4129 ( n8327 , n5574 );
    not g4130 ( n14236 , n28285 );
    not g4131 ( n27856 , n17117 );
    not g4132 ( n11049 , n11800 );
    and g4133 ( n25479 , n24405 , n16338 );
    not g4134 ( n18941 , n1670 );
    or g4135 ( n26868 , n13821 , n21732 );
    or g4136 ( n13056 , n22331 , n16123 );
    xor g4137 ( n4089 , n17759 , n24429 );
    or g4138 ( n16102 , n22624 , n2399 );
    xnor g4139 ( n269 , n30103 , n23851 );
    and g4140 ( n15412 , n16669 , n27341 );
    and g4141 ( n9186 , n14759 , n28669 );
    xor g4142 ( n20714 , n4427 , n27386 );
    and g4143 ( n989 , n7442 , n20151 );
    xnor g4144 ( n5581 , n4392 , n19853 );
    nor g4145 ( n15069 , n4554 , n25982 );
    or g4146 ( n21219 , n31384 , n25823 );
    and g4147 ( n14969 , n9198 , n27174 );
    xnor g4148 ( n30564 , n20957 , n10413 );
    not g4149 ( n29728 , n4594 );
    not g4150 ( n9960 , n10479 );
    or g4151 ( n5151 , n1285 , n10236 );
    xnor g4152 ( n24891 , n18781 , n18986 );
    not g4153 ( n21551 , n20155 );
    not g4154 ( n427 , n20431 );
    or g4155 ( n7498 , n7295 , n1766 );
    xnor g4156 ( n12259 , n9602 , n14695 );
    or g4157 ( n12931 , n30706 , n13859 );
    or g4158 ( n12334 , n9655 , n30934 );
    not g4159 ( n6737 , n25883 );
    not g4160 ( n3870 , n7087 );
    and g4161 ( n15008 , n25400 , n28187 );
    xnor g4162 ( n21726 , n17944 , n25469 );
    xnor g4163 ( n31156 , n3061 , n4951 );
    and g4164 ( n24372 , n7412 , n22857 );
    and g4165 ( n16534 , n4204 , n31333 );
    and g4166 ( n15440 , n19195 , n11895 );
    or g4167 ( n8741 , n7354 , n8867 );
    or g4168 ( n13722 , n23561 , n12879 );
    not g4169 ( n7794 , n14547 );
    or g4170 ( n6363 , n30227 , n2089 );
    or g4171 ( n10583 , n3953 , n7499 );
    xnor g4172 ( n21867 , n8008 , n29363 );
    not g4173 ( n17018 , n13029 );
    not g4174 ( n9276 , n29444 );
    not g4175 ( n4204 , n10483 );
    or g4176 ( n13253 , n28512 , n30021 );
    and g4177 ( n4671 , n19451 , n809 );
    or g4178 ( n1503 , n19330 , n11474 );
    nor g4179 ( n20373 , n13635 , n30546 );
    xnor g4180 ( n26413 , n14922 , n189 );
    and g4181 ( n6664 , n19991 , n5342 );
    or g4182 ( n10089 , n28428 , n17077 );
    or g4183 ( n20980 , n4141 , n22247 );
    or g4184 ( n16378 , n6282 , n29362 );
    xnor g4185 ( n28845 , n25896 , n12607 );
    and g4186 ( n1289 , n26045 , n28728 );
    or g4187 ( n31632 , n24040 , n26917 );
    nor g4188 ( n19426 , n24246 , n11574 );
    not g4189 ( n13188 , n30720 );
    and g4190 ( n7096 , n12175 , n30201 );
    or g4191 ( n6631 , n7385 , n24087 );
    xnor g4192 ( n23375 , n25139 , n30989 );
    not g4193 ( n12133 , n18201 );
    not g4194 ( n26163 , n5006 );
    or g4195 ( n79 , n6873 , n29629 );
    not g4196 ( n11250 , n30894 );
    buf g4197 ( n16193 , n2058 );
    xnor g4198 ( n16205 , n25856 , n25793 );
    xnor g4199 ( n4292 , n11658 , n28006 );
    or g4200 ( n20257 , n4519 , n7681 );
    not g4201 ( n21131 , n25577 );
    nor g4202 ( n13373 , n29389 , n9620 );
    not g4203 ( n26523 , n23681 );
    not g4204 ( n5870 , n28843 );
    not g4205 ( n11069 , n14474 );
    not g4206 ( n9417 , n16189 );
    or g4207 ( n22898 , n15598 , n24630 );
    or g4208 ( n9649 , n25441 , n25376 );
    xnor g4209 ( n20832 , n6229 , n16270 );
    not g4210 ( n13283 , n28095 );
    nor g4211 ( n24384 , n24129 , n7930 );
    xnor g4212 ( n27569 , n4157 , n5792 );
    and g4213 ( n13106 , n3651 , n18930 );
    or g4214 ( n9308 , n15588 , n8403 );
    xnor g4215 ( n31573 , n2618 , n9970 );
    xnor g4216 ( n7093 , n7103 , n3269 );
    and g4217 ( n30582 , n7305 , n10448 );
    xor g4218 ( n1678 , n20817 , n7875 );
    and g4219 ( n22003 , n31776 , n24374 );
    nor g4220 ( n19048 , n13573 , n20659 );
    or g4221 ( n19403 , n29033 , n20634 );
    xor g4222 ( n18735 , n931 , n614 );
    xnor g4223 ( n19170 , n19516 , n7046 );
    not g4224 ( n13172 , n6306 );
    or g4225 ( n19387 , n31832 , n7257 );
    xnor g4226 ( n19428 , n16639 , n12409 );
    xnor g4227 ( n14589 , n3399 , n29524 );
    not g4228 ( n27250 , n14356 );
    or g4229 ( n26892 , n10059 , n19816 );
    or g4230 ( n23011 , n2483 , n946 );
    or g4231 ( n4167 , n2119 , n24713 );
    xnor g4232 ( n19460 , n27418 , n7766 );
    not g4233 ( n27204 , n24871 );
    and g4234 ( n27634 , n24469 , n12161 );
    not g4235 ( n14026 , n13137 );
    nor g4236 ( n4164 , n5406 , n1774 );
    and g4237 ( n24337 , n22426 , n26697 );
    or g4238 ( n26692 , n5338 , n13174 );
    xnor g4239 ( n21370 , n18357 , n3649 );
    nor g4240 ( n11235 , n20913 , n16041 );
    or g4241 ( n11310 , n4232 , n28540 );
    xnor g4242 ( n22849 , n18388 , n30685 );
    not g4243 ( n25497 , n9684 );
    and g4244 ( n14990 , n10170 , n26739 );
    or g4245 ( n6417 , n31060 , n13300 );
    and g4246 ( n22861 , n2979 , n6116 );
    buf g4247 ( n11850 , n25596 );
    not g4248 ( n13616 , n12806 );
    xnor g4249 ( n26939 , n26004 , n30411 );
    xnor g4250 ( n11025 , n29941 , n3653 );
    not g4251 ( n29493 , n29073 );
    or g4252 ( n29579 , n3679 , n1075 );
    not g4253 ( n9706 , n11139 );
    not g4254 ( n28372 , n1433 );
    or g4255 ( n22949 , n19668 , n4614 );
    and g4256 ( n6524 , n4372 , n15108 );
    xnor g4257 ( n21490 , n26002 , n1095 );
    buf g4258 ( n3059 , n31353 );
    nor g4259 ( n12544 , n30604 , n27864 );
    xnor g4260 ( n5231 , n22951 , n7282 );
    and g4261 ( n10796 , n10606 , n23001 );
    or g4262 ( n12714 , n12668 , n27086 );
    not g4263 ( n31851 , n27233 );
    or g4264 ( n24390 , n30312 , n5769 );
    nor g4265 ( n29921 , n8664 , n22820 );
    not g4266 ( n4216 , n10321 );
    not g4267 ( n27947 , n14184 );
    not g4268 ( n12593 , n28791 );
    and g4269 ( n11786 , n16102 , n22513 );
    buf g4270 ( n12318 , n27818 );
    or g4271 ( n19528 , n20621 , n3305 );
    and g4272 ( n24413 , n25011 , n24783 );
    and g4273 ( n12537 , n4167 , n19052 );
    not g4274 ( n10508 , n11743 );
    not g4275 ( n2395 , n2963 );
    xnor g4276 ( n29212 , n27911 , n3475 );
    not g4277 ( n18447 , n8540 );
    xnor g4278 ( n31654 , n11028 , n17305 );
    not g4279 ( n4804 , n5418 );
    xnor g4280 ( n6736 , n3848 , n31709 );
    or g4281 ( n10012 , n11728 , n23875 );
    or g4282 ( n970 , n27885 , n26996 );
    and g4283 ( n15430 , n18481 , n14023 );
    or g4284 ( n4062 , n7663 , n14100 );
    not g4285 ( n29335 , n18485 );
    or g4286 ( n27220 , n12710 , n24420 );
    or g4287 ( n24424 , n31259 , n4067 );
    or g4288 ( n7615 , n4869 , n17315 );
    or g4289 ( n19442 , n6108 , n18945 );
    or g4290 ( n9921 , n23887 , n10175 );
    or g4291 ( n22289 , n8603 , n13177 );
    nor g4292 ( n22474 , n30908 , n7692 );
    not g4293 ( n20485 , n14815 );
    or g4294 ( n5020 , n23259 , n24166 );
    not g4295 ( n16273 , n7351 );
    or g4296 ( n24731 , n20826 , n11820 );
    not g4297 ( n8084 , n31416 );
    xnor g4298 ( n28720 , n19626 , n24272 );
    not g4299 ( n1378 , n23789 );
    and g4300 ( n12894 , n10663 , n6812 );
    and g4301 ( n14222 , n3464 , n5313 );
    or g4302 ( n17635 , n15638 , n29241 );
    and g4303 ( n30133 , n23497 , n25897 );
    or g4304 ( n13525 , n10787 , n9506 );
    nor g4305 ( n25325 , n14361 , n26769 );
    or g4306 ( n30017 , n7531 , n14394 );
    or g4307 ( n6785 , n8037 , n12028 );
    or g4308 ( n18630 , n30881 , n26278 );
    or g4309 ( n21715 , n26612 , n26195 );
    not g4310 ( n22503 , n24213 );
    and g4311 ( n9256 , n22062 , n10280 );
    not g4312 ( n7525 , n6535 );
    and g4313 ( n29035 , n6887 , n13173 );
    or g4314 ( n13783 , n29818 , n10630 );
    or g4315 ( n11616 , n12024 , n23900 );
    and g4316 ( n641 , n10192 , n19972 );
    and g4317 ( n25906 , n18030 , n18316 );
    or g4318 ( n8643 , n6006 , n6615 );
    not g4319 ( n7958 , n29 );
    or g4320 ( n13652 , n20887 , n14126 );
    and g4321 ( n29160 , n5154 , n8098 );
    and g4322 ( n9284 , n14889 , n19199 );
    xnor g4323 ( n30431 , n26799 , n31671 );
    xnor g4324 ( n1744 , n13819 , n23759 );
    not g4325 ( n28315 , n3698 );
    or g4326 ( n4826 , n29688 , n31350 );
    and g4327 ( n29408 , n4537 , n19169 );
    xnor g4328 ( n2608 , n31585 , n6331 );
    and g4329 ( n2955 , n29456 , n8107 );
    or g4330 ( n10087 , n6271 , n7222 );
    or g4331 ( n25357 , n12095 , n29773 );
    nor g4332 ( n8482 , n31474 , n12184 );
    or g4333 ( n23238 , n30024 , n14765 );
    not g4334 ( n14823 , n12087 );
    not g4335 ( n8553 , n7592 );
    xnor g4336 ( n416 , n30438 , n1860 );
    and g4337 ( n3327 , n31488 , n26022 );
    not g4338 ( n642 , n29153 );
    xnor g4339 ( n30351 , n29444 , n7314 );
    or g4340 ( n5537 , n31226 , n6380 );
    and g4341 ( n5830 , n31011 , n25723 );
    xnor g4342 ( n13277 , n29172 , n16815 );
    xnor g4343 ( n16587 , n14607 , n30590 );
    nor g4344 ( n10070 , n1177 , n7274 );
    or g4345 ( n28358 , n20630 , n2160 );
    not g4346 ( n20482 , n6511 );
    not g4347 ( n8712 , n31970 );
    not g4348 ( n26916 , n17811 );
    nor g4349 ( n3292 , n21105 , n19502 );
    xor g4350 ( n29117 , n28136 , n1177 );
    not g4351 ( n13987 , n12993 );
    nor g4352 ( n7543 , n31725 , n18385 );
    nor g4353 ( n17852 , n16029 , n8360 );
    or g4354 ( n6897 , n1372 , n16087 );
    and g4355 ( n31192 , n19101 , n18388 );
    xnor g4356 ( n18829 , n11941 , n571 );
    nor g4357 ( n13350 , n28267 , n17896 );
    or g4358 ( n17247 , n14509 , n10224 );
    or g4359 ( n15042 , n225 , n24170 );
    or g4360 ( n15565 , n2849 , n30975 );
    and g4361 ( n14592 , n15371 , n4753 );
    or g4362 ( n7590 , n6959 , n16371 );
    xnor g4363 ( n4391 , n6678 , n29310 );
    not g4364 ( n7877 , n8284 );
    nor g4365 ( n13484 , n30674 , n1 );
    xnor g4366 ( n7513 , n21153 , n15500 );
    xnor g4367 ( n26812 , n18721 , n12153 );
    xnor g4368 ( n7101 , n29245 , n29066 );
    not g4369 ( n27609 , n17847 );
    not g4370 ( n13111 , n26486 );
    or g4371 ( n15294 , n14192 , n602 );
    or g4372 ( n10819 , n8870 , n22087 );
    xnor g4373 ( n24349 , n24455 , n21708 );
    buf g4374 ( n23423 , n11187 );
    nor g4375 ( n18649 , n31731 , n1375 );
    xor g4376 ( n16125 , n16827 , n7965 );
    not g4377 ( n9528 , n6342 );
    xnor g4378 ( n25883 , n8277 , n5256 );
    nor g4379 ( n147 , n21075 , n8644 );
    nor g4380 ( n4163 , n9889 , n10228 );
    and g4381 ( n26404 , n19114 , n12888 );
    not g4382 ( n31155 , n28977 );
    not g4383 ( n25072 , n3755 );
    xnor g4384 ( n29304 , n15573 , n1973 );
    xnor g4385 ( n28783 , n23687 , n11137 );
    not g4386 ( n16126 , n9195 );
    xnor g4387 ( n17633 , n18551 , n23306 );
    not g4388 ( n17125 , n31160 );
    or g4389 ( n517 , n21462 , n17626 );
    or g4390 ( n24352 , n4372 , n13493 );
    not g4391 ( n23638 , n18920 );
    not g4392 ( n8114 , n20071 );
    buf g4393 ( n22841 , n8824 );
    or g4394 ( n14628 , n18241 , n15364 );
    xnor g4395 ( n22677 , n14069 , n14828 );
    not g4396 ( n30934 , n12030 );
    or g4397 ( n23506 , n15506 , n3985 );
    nor g4398 ( n28254 , n8014 , n8514 );
    and g4399 ( n10264 , n7294 , n2215 );
    not g4400 ( n29635 , n28937 );
    or g4401 ( n8170 , n8716 , n9457 );
    or g4402 ( n14101 , n10290 , n14645 );
    xnor g4403 ( n31854 , n19750 , n23615 );
    xnor g4404 ( n12686 , n4415 , n14203 );
    buf g4405 ( n717 , n29192 );
    and g4406 ( n16571 , n3043 , n14711 );
    xnor g4407 ( n17805 , n26843 , n25378 );
    or g4408 ( n22317 , n29517 , n14494 );
    nor g4409 ( n23090 , n11438 , n7661 );
    or g4410 ( n21651 , n11886 , n27250 );
    xnor g4411 ( n3800 , n4591 , n25200 );
    nor g4412 ( n11314 , n25305 , n14523 );
    not g4413 ( n4115 , n26460 );
    xnor g4414 ( n26301 , n31411 , n469 );
    xnor g4415 ( n31661 , n3284 , n14373 );
    and g4416 ( n30438 , n1649 , n12740 );
    not g4417 ( n23723 , n17213 );
    xnor g4418 ( n25311 , n28829 , n862 );
    or g4419 ( n19828 , n2010 , n19683 );
    or g4420 ( n3325 , n6452 , n8022 );
    xnor g4421 ( n31313 , n14879 , n25197 );
    nor g4422 ( n13334 , n793 , n8440 );
    xnor g4423 ( n8592 , n8036 , n31380 );
    or g4424 ( n16743 , n2017 , n30898 );
    not g4425 ( n14585 , n28804 );
    buf g4426 ( n344 , n12725 );
    or g4427 ( n2172 , n31616 , n3546 );
    not g4428 ( n19928 , n21588 );
    xnor g4429 ( n14796 , n8951 , n10232 );
    xnor g4430 ( n1946 , n26763 , n7414 );
    or g4431 ( n29983 , n3271 , n21430 );
    not g4432 ( n26428 , n26306 );
    or g4433 ( n4553 , n24118 , n23954 );
    not g4434 ( n4809 , n27256 );
    not g4435 ( n3428 , n19891 );
    not g4436 ( n5989 , n7796 );
    not g4437 ( n14083 , n29290 );
    or g4438 ( n9722 , n22838 , n23301 );
    not g4439 ( n936 , n10269 );
    or g4440 ( n10587 , n9802 , n18358 );
    or g4441 ( n27294 , n19439 , n19531 );
    not g4442 ( n30036 , n3587 );
    and g4443 ( n20072 , n17643 , n21082 );
    or g4444 ( n31312 , n15894 , n7517 );
    xnor g4445 ( n1709 , n9168 , n17867 );
    not g4446 ( n25531 , n29307 );
    xnor g4447 ( n591 , n27735 , n2091 );
    or g4448 ( n24580 , n23358 , n16953 );
    not g4449 ( n8907 , n2064 );
    not g4450 ( n19732 , n13759 );
    or g4451 ( n10143 , n15625 , n330 );
    and g4452 ( n6293 , n7406 , n23517 );
    nor g4453 ( n5016 , n6127 , n8407 );
    not g4454 ( n28486 , n5375 );
    or g4455 ( n22531 , n26330 , n732 );
    xnor g4456 ( n9554 , n23466 , n22901 );
    nor g4457 ( n9567 , n16131 , n26487 );
    not g4458 ( n14011 , n3350 );
    or g4459 ( n22407 , n22744 , n17693 );
    or g4460 ( n27353 , n30177 , n4841 );
    not g4461 ( n16839 , n9321 );
    xnor g4462 ( n5230 , n8098 , n29702 );
    or g4463 ( n18390 , n3296 , n9271 );
    xnor g4464 ( n29968 , n9417 , n22886 );
    and g4465 ( n3134 , n13249 , n31826 );
    not g4466 ( n28818 , n6226 );
    and g4467 ( n27745 , n25651 , n19792 );
    or g4468 ( n12386 , n5720 , n13596 );
    not g4469 ( n4653 , n16413 );
    nor g4470 ( n27810 , n16315 , n19034 );
    nor g4471 ( n23563 , n20790 , n18373 );
    or g4472 ( n1822 , n13872 , n11620 );
    or g4473 ( n22177 , n16374 , n277 );
    nor g4474 ( n26236 , n3641 , n3033 );
    not g4475 ( n15803 , n6826 );
    or g4476 ( n5513 , n31553 , n31068 );
    xnor g4477 ( n31415 , n25777 , n3293 );
    xnor g4478 ( n17224 , n15588 , n13700 );
    xor g4479 ( n14328 , n22112 , n238 );
    and g4480 ( n16114 , n27995 , n9773 );
    not g4481 ( n12773 , n29919 );
    and g4482 ( n2332 , n30580 , n10098 );
    not g4483 ( n31901 , n988 );
    xnor g4484 ( n27748 , n20482 , n9743 );
    xnor g4485 ( n8508 , n20859 , n13888 );
    not g4486 ( n11816 , n29426 );
    not g4487 ( n12961 , n19516 );
    or g4488 ( n21331 , n10765 , n24085 );
    or g4489 ( n23445 , n7568 , n21948 );
    nor g4490 ( n4850 , n22355 , n26391 );
    xnor g4491 ( n17526 , n28370 , n2444 );
    not g4492 ( n8948 , n21192 );
    xnor g4493 ( n5481 , n2932 , n10781 );
    and g4494 ( n10419 , n26397 , n24193 );
    or g4495 ( n30755 , n16230 , n10085 );
    xnor g4496 ( n31937 , n24118 , n28734 );
    or g4497 ( n2651 , n1069 , n9413 );
    not g4498 ( n1532 , n29393 );
    xnor g4499 ( n19352 , n17432 , n19425 );
    xnor g4500 ( n28269 , n26040 , n15453 );
    and g4501 ( n16121 , n2140 , n25005 );
    and g4502 ( n26088 , n17076 , n10493 );
    or g4503 ( n9521 , n11425 , n19701 );
    nor g4504 ( n7870 , n16730 , n9200 );
    or g4505 ( n23030 , n30807 , n20671 );
    and g4506 ( n12721 , n23775 , n3090 );
    or g4507 ( n15879 , n7104 , n9367 );
    not g4508 ( n9475 , n11512 );
    and g4509 ( n4244 , n8027 , n29105 );
    xnor g4510 ( n21021 , n22188 , n27510 );
    not g4511 ( n5525 , n24104 );
    not g4512 ( n21264 , n21849 );
    or g4513 ( n30450 , n10309 , n22400 );
    not g4514 ( n4803 , n18886 );
    xnor g4515 ( n30753 , n4275 , n29553 );
    xnor g4516 ( n19755 , n12041 , n14842 );
    not g4517 ( n14763 , n12951 );
    not g4518 ( n16000 , n11609 );
    and g4519 ( n5769 , n8206 , n14849 );
    not g4520 ( n7159 , n13073 );
    not g4521 ( n28637 , n2255 );
    nor g4522 ( n21143 , n9324 , n21551 );
    not g4523 ( n13534 , n5299 );
    or g4524 ( n16497 , n27243 , n25154 );
    and g4525 ( n3586 , n14009 , n24126 );
    not g4526 ( n28973 , n14657 );
    not g4527 ( n19042 , n27126 );
    xnor g4528 ( n5062 , n27640 , n18444 );
    or g4529 ( n19839 , n16276 , n22491 );
    and g4530 ( n15177 , n11615 , n25894 );
    not g4531 ( n18202 , n23852 );
    and g4532 ( n1133 , n7627 , n31341 );
    and g4533 ( n1438 , n9296 , n17562 );
    or g4534 ( n25617 , n7026 , n6254 );
    or g4535 ( n7869 , n28880 , n20288 );
    not g4536 ( n10664 , n20804 );
    not g4537 ( n16424 , n27155 );
    xnor g4538 ( n30404 , n29444 , n24794 );
    and g4539 ( n1108 , n19653 , n26199 );
    not g4540 ( n3355 , n25165 );
    and g4541 ( n17377 , n360 , n24597 );
    and g4542 ( n28175 , n19799 , n16244 );
    not g4543 ( n6947 , n24909 );
    and g4544 ( n569 , n29624 , n2909 );
    not g4545 ( n1143 , n17758 );
    or g4546 ( n12257 , n11967 , n4268 );
    xor g4547 ( n1231 , n25778 , n31535 );
    or g4548 ( n23004 , n10060 , n12151 );
    or g4549 ( n12785 , n28341 , n29866 );
    and g4550 ( n8271 , n25440 , n18894 );
    or g4551 ( n10023 , n18055 , n20389 );
    or g4552 ( n12966 , n25334 , n1006 );
    and g4553 ( n16819 , n12354 , n24889 );
    and g4554 ( n9393 , n6992 , n18443 );
    and g4555 ( n13738 , n15414 , n10731 );
    or g4556 ( n22888 , n29353 , n17192 );
    nor g4557 ( n14719 , n16182 , n289 );
    not g4558 ( n12649 , n23724 );
    xnor g4559 ( n18926 , n18122 , n19911 );
    xnor g4560 ( n24113 , n16513 , n15927 );
    xnor g4561 ( n7931 , n27676 , n24947 );
    or g4562 ( n20537 , n10503 , n136 );
    and g4563 ( n7144 , n8864 , n16588 );
    not g4564 ( n18357 , n25164 );
    not g4565 ( n29356 , n22418 );
    or g4566 ( n19971 , n21235 , n28323 );
    or g4567 ( n1617 , n7859 , n5895 );
    not g4568 ( n31062 , n2447 );
    not g4569 ( n27549 , n9011 );
    not g4570 ( n26889 , n28712 );
    and g4571 ( n8015 , n7612 , n30480 );
    xnor g4572 ( n7857 , n20879 , n27836 );
    not g4573 ( n1869 , n18331 );
    xnor g4574 ( n19731 , n6061 , n28417 );
    xnor g4575 ( n4711 , n171 , n23732 );
    xnor g4576 ( n14774 , n14372 , n27481 );
    xnor g4577 ( n2569 , n19381 , n27010 );
    not g4578 ( n29426 , n21923 );
    xnor g4579 ( n17336 , n27716 , n8804 );
    and g4580 ( n28129 , n4043 , n701 );
    not g4581 ( n5246 , n25035 );
    or g4582 ( n4438 , n5363 , n24673 );
    or g4583 ( n31599 , n17710 , n10855 );
    or g4584 ( n31587 , n9338 , n14362 );
    xnor g4585 ( n8469 , n18881 , n8030 );
    xnor g4586 ( n7291 , n13325 , n11054 );
    xnor g4587 ( n18734 , n13288 , n4987 );
    xnor g4588 ( n30543 , n26046 , n9477 );
    xnor g4589 ( n2388 , n10822 , n7387 );
    and g4590 ( n9413 , n6017 , n28996 );
    xnor g4591 ( n31881 , n6740 , n18914 );
    xnor g4592 ( n27847 , n23360 , n6098 );
    or g4593 ( n20415 , n30514 , n24510 );
    not g4594 ( n11393 , n27275 );
    xnor g4595 ( n16387 , n18717 , n23489 );
    nor g4596 ( n28249 , n28004 , n29766 );
    nor g4597 ( n21930 , n8919 , n2372 );
    xnor g4598 ( n11177 , n24623 , n1961 );
    or g4599 ( n21194 , n13669 , n5786 );
    or g4600 ( n13442 , n23825 , n62 );
    and g4601 ( n4852 , n15850 , n22703 );
    nor g4602 ( n11489 , n16805 , n9621 );
    not g4603 ( n11704 , n21726 );
    xnor g4604 ( n27721 , n14503 , n20365 );
    xnor g4605 ( n17705 , n24630 , n1039 );
    not g4606 ( n17102 , n3361 );
    or g4607 ( n20550 , n1011 , n1598 );
    not g4608 ( n11259 , n12680 );
    not g4609 ( n18643 , n1427 );
    xnor g4610 ( n10899 , n1886 , n16973 );
    and g4611 ( n11879 , n2279 , n7826 );
    not g4612 ( n31678 , n6904 );
    or g4613 ( n23592 , n9428 , n29255 );
    nor g4614 ( n1431 , n17910 , n21384 );
    not g4615 ( n25104 , n24624 );
    or g4616 ( n31766 , n1150 , n16727 );
    or g4617 ( n16816 , n16026 , n15279 );
    and g4618 ( n18085 , n24142 , n27111 );
    and g4619 ( n29860 , n6753 , n13460 );
    not g4620 ( n6689 , n15024 );
    xnor g4621 ( n26524 , n16453 , n2836 );
    nor g4622 ( n1721 , n4723 , n21297 );
    xnor g4623 ( n29580 , n27233 , n12777 );
    not g4624 ( n21646 , n18362 );
    or g4625 ( n6656 , n19612 , n11910 );
    xnor g4626 ( n3121 , n31992 , n12627 );
    or g4627 ( n24256 , n20177 , n1530 );
    not g4628 ( n2524 , n25028 );
    not g4629 ( n9716 , n14841 );
    and g4630 ( n24815 , n2865 , n30626 );
    and g4631 ( n3788 , n16120 , n6238 );
    and g4632 ( n29135 , n22329 , n18872 );
    or g4633 ( n7203 , n26438 , n28385 );
    not g4634 ( n21671 , n14670 );
    and g4635 ( n28853 , n1085 , n245 );
    xnor g4636 ( n26860 , n9939 , n12072 );
    not g4637 ( n19406 , n1430 );
    xnor g4638 ( n8433 , n27552 , n22547 );
    not g4639 ( n30690 , n29967 );
    and g4640 ( n28814 , n3507 , n1657 );
    nor g4641 ( n8565 , n23419 , n17289 );
    not g4642 ( n12383 , n13594 );
    nor g4643 ( n17143 , n23223 , n11899 );
    and g4644 ( n11072 , n10432 , n31500 );
    and g4645 ( n30751 , n22195 , n30736 );
    and g4646 ( n20783 , n25737 , n12206 );
    or g4647 ( n9340 , n25285 , n148 );
    xnor g4648 ( n30941 , n8680 , n16454 );
    xnor g4649 ( n12546 , n16347 , n19221 );
    and g4650 ( n20497 , n8145 , n18057 );
    nor g4651 ( n26326 , n15382 , n17032 );
    xor g4652 ( n7351 , n9343 , n28137 );
    not g4653 ( n11389 , n2858 );
    and g4654 ( n25957 , n21495 , n1965 );
    xnor g4655 ( n1066 , n24979 , n22798 );
    and g4656 ( n1498 , n13989 , n13536 );
    xnor g4657 ( n10365 , n19499 , n24244 );
    not g4658 ( n12677 , n202 );
    and g4659 ( n4877 , n12381 , n31658 );
    or g4660 ( n1155 , n13109 , n5129 );
    or g4661 ( n13571 , n31511 , n24649 );
    not g4662 ( n3885 , n311 );
    nor g4663 ( n19246 , n21679 , n7104 );
    not g4664 ( n4755 , n10611 );
    xnor g4665 ( n27868 , n15480 , n1810 );
    and g4666 ( n25606 , n25901 , n24373 );
    xnor g4667 ( n8081 , n31899 , n16100 );
    xnor g4668 ( n26385 , n6071 , n6145 );
    not g4669 ( n26445 , n21003 );
    not g4670 ( n2049 , n6957 );
    xnor g4671 ( n28135 , n8073 , n23798 );
    xnor g4672 ( n5334 , n26413 , n9591 );
    and g4673 ( n23014 , n27865 , n8561 );
    and g4674 ( n24670 , n14848 , n25552 );
    or g4675 ( n23665 , n28329 , n31084 );
    nor g4676 ( n19308 , n9310 , n10737 );
    xnor g4677 ( n7387 , n4895 , n2898 );
    or g4678 ( n830 , n17149 , n18001 );
    xnor g4679 ( n26121 , n10465 , n8400 );
    not g4680 ( n2617 , n9540 );
    and g4681 ( n30137 , n8962 , n28650 );
    or g4682 ( n30307 , n6634 , n1379 );
    or g4683 ( n16145 , n30882 , n13512 );
    xnor g4684 ( n31105 , n9881 , n8808 );
    and g4685 ( n25442 , n7738 , n19571 );
    or g4686 ( n4965 , n18434 , n27585 );
    not g4687 ( n13448 , n31327 );
    or g4688 ( n8303 , n15880 , n2761 );
    not g4689 ( n12533 , n27318 );
    or g4690 ( n2413 , n5594 , n24002 );
    or g4691 ( n4801 , n25957 , n17707 );
    nor g4692 ( n16537 , n3755 , n28260 );
    not g4693 ( n13475 , n9362 );
    xnor g4694 ( n26530 , n5740 , n30311 );
    or g4695 ( n22062 , n29315 , n3180 );
    not g4696 ( n7983 , n31548 );
    or g4697 ( n11009 , n27077 , n12728 );
    and g4698 ( n16569 , n11993 , n28293 );
    not g4699 ( n993 , n24520 );
    or g4700 ( n22414 , n31797 , n23202 );
    or g4701 ( n484 , n5251 , n9809 );
    nor g4702 ( n6586 , n19182 , n12609 );
    not g4703 ( n20165 , n4125 );
    not g4704 ( n24306 , n15687 );
    not g4705 ( n6594 , n5276 );
    and g4706 ( n21360 , n13115 , n15188 );
    or g4707 ( n4506 , n15940 , n2287 );
    not g4708 ( n3288 , n7369 );
    or g4709 ( n8590 , n19071 , n6097 );
    nor g4710 ( n12330 , n14133 , n18246 );
    and g4711 ( n10186 , n18073 , n12957 );
    or g4712 ( n43 , n10430 , n30444 );
    xnor g4713 ( n15869 , n13210 , n20181 );
    and g4714 ( n27700 , n17463 , n7976 );
    xnor g4715 ( n3022 , n21848 , n13277 );
    not g4716 ( n19871 , n31853 );
    nor g4717 ( n9204 , n12888 , n21819 );
    not g4718 ( n14089 , n22802 );
    xnor g4719 ( n8510 , n28716 , n20096 );
    xnor g4720 ( n28045 , n16856 , n3996 );
    not g4721 ( n526 , n14225 );
    not g4722 ( n21375 , n4749 );
    not g4723 ( n12919 , n12758 );
    not g4724 ( n24894 , n25006 );
    and g4725 ( n1239 , n22540 , n22008 );
    not g4726 ( n18329 , n6260 );
    not g4727 ( n254 , n13321 );
    or g4728 ( n29222 , n16197 , n23525 );
    or g4729 ( n5802 , n16215 , n14382 );
    xnor g4730 ( n23148 , n9591 , n3688 );
    not g4731 ( n21598 , n20029 );
    xnor g4732 ( n4453 , n21374 , n27538 );
    not g4733 ( n28242 , n13495 );
    and g4734 ( n17288 , n11364 , n15302 );
    or g4735 ( n12548 , n23010 , n29926 );
    xor g4736 ( n30426 , n7335 , n13902 );
    nor g4737 ( n11258 , n24578 , n21134 );
    xnor g4738 ( n5758 , n4363 , n12076 );
    nor g4739 ( n6855 , n25654 , n16564 );
    not g4740 ( n4071 , n10470 );
    and g4741 ( n3343 , n18111 , n19685 );
    xor g4742 ( n29785 , n6255 , n13760 );
    xnor g4743 ( n4935 , n19836 , n18570 );
    not g4744 ( n4628 , n29196 );
    not g4745 ( n23169 , n614 );
    xnor g4746 ( n3400 , n3758 , n19471 );
    not g4747 ( n18255 , n11636 );
    xnor g4748 ( n7849 , n18373 , n11711 );
    not g4749 ( n25103 , n18504 );
    or g4750 ( n17609 , n7764 , n24041 );
    xnor g4751 ( n6298 , n17825 , n5192 );
    nor g4752 ( n20995 , n8397 , n9674 );
    or g4753 ( n29858 , n13359 , n21157 );
    xnor g4754 ( n19891 , n13804 , n22315 );
    xor g4755 ( n13843 , n16000 , n18850 );
    or g4756 ( n31378 , n16236 , n26761 );
    not g4757 ( n25372 , n21914 );
    or g4758 ( n28733 , n12625 , n4619 );
    or g4759 ( n29174 , n30096 , n1020 );
    xnor g4760 ( n25453 , n2830 , n5812 );
    not g4761 ( n1347 , n7692 );
    not g4762 ( n13539 , n27448 );
    xnor g4763 ( n12425 , n22839 , n15207 );
    xnor g4764 ( n22577 , n7556 , n778 );
    not g4765 ( n31382 , n23549 );
    or g4766 ( n5584 , n27318 , n9527 );
    not g4767 ( n13192 , n16563 );
    or g4768 ( n10578 , n6041 , n21562 );
    or g4769 ( n27059 , n12184 , n23912 );
    xnor g4770 ( n30837 , n21198 , n28497 );
    or g4771 ( n5195 , n13701 , n26070 );
    xnor g4772 ( n21191 , n8386 , n13765 );
    or g4773 ( n17562 , n23852 , n14290 );
    and g4774 ( n6913 , n23977 , n2661 );
    xnor g4775 ( n10120 , n17237 , n4239 );
    or g4776 ( n20228 , n6331 , n2606 );
    not g4777 ( n8540 , n13814 );
    xnor g4778 ( n7113 , n22917 , n3345 );
    or g4779 ( n10646 , n21428 , n5983 );
    or g4780 ( n26680 , n17567 , n16641 );
    not g4781 ( n24165 , n17601 );
    not g4782 ( n14155 , n9202 );
    and g4783 ( n15963 , n16388 , n9128 );
    nor g4784 ( n4060 , n7335 , n2640 );
    xnor g4785 ( n16068 , n20377 , n29458 );
    not g4786 ( n28864 , n1018 );
    or g4787 ( n19515 , n3637 , n26611 );
    xnor g4788 ( n29318 , n28755 , n16815 );
    or g4789 ( n14207 , n29999 , n23721 );
    or g4790 ( n6663 , n21314 , n14507 );
    not g4791 ( n21712 , n26658 );
    not g4792 ( n6650 , n20795 );
    and g4793 ( n15961 , n18188 , n5497 );
    or g4794 ( n21498 , n20967 , n21726 );
    or g4795 ( n28664 , n23677 , n28927 );
    xor g4796 ( n144 , n19915 , n14653 );
    xnor g4797 ( n19562 , n10363 , n14711 );
    xnor g4798 ( n21903 , n20837 , n18725 );
    or g4799 ( n19037 , n282 , n2686 );
    xnor g4800 ( n3619 , n13467 , n25579 );
    not g4801 ( n23297 , n7974 );
    xnor g4802 ( n16359 , n14598 , n27368 );
    xor g4803 ( n15733 , n14139 , n21418 );
    or g4804 ( n5961 , n4016 , n27703 );
    xnor g4805 ( n11519 , n25854 , n14945 );
    nor g4806 ( n31292 , n26004 , n22497 );
    and g4807 ( n10541 , n17810 , n18745 );
    nor g4808 ( n17997 , n11792 , n12564 );
    not g4809 ( n8973 , n4251 );
    or g4810 ( n23589 , n17851 , n25239 );
    or g4811 ( n16606 , n28248 , n9084 );
    not g4812 ( n22073 , n22641 );
    or g4813 ( n2730 , n25979 , n1311 );
    or g4814 ( n25944 , n7120 , n19259 );
    xnor g4815 ( n2100 , n29154 , n15012 );
    nor g4816 ( n18687 , n20080 , n28 );
    not g4817 ( n11504 , n21249 );
    not g4818 ( n327 , n21058 );
    xnor g4819 ( n27517 , n1195 , n3163 );
    and g4820 ( n22333 , n18556 , n10995 );
    xor g4821 ( n23639 , n29354 , n21096 );
    not g4822 ( n9986 , n9354 );
    xnor g4823 ( n6112 , n7904 , n238 );
    not g4824 ( n11976 , n24596 );
    xnor g4825 ( n26626 , n64 , n25276 );
    not g4826 ( n15122 , n20526 );
    not g4827 ( n7839 , n25257 );
    not g4828 ( n29476 , n30575 );
    not g4829 ( n26976 , n7447 );
    xnor g4830 ( n2864 , n3496 , n26814 );
    xnor g4831 ( n10687 , n19615 , n31481 );
    xor g4832 ( n18385 , n16257 , n31593 );
    not g4833 ( n18396 , n17862 );
    or g4834 ( n28972 , n14474 , n11595 );
    xnor g4835 ( n9118 , n2468 , n4547 );
    not g4836 ( n26353 , n7077 );
    xnor g4837 ( n18658 , n25598 , n31690 );
    and g4838 ( n23062 , n22915 , n15321 );
    xnor g4839 ( n9588 , n25463 , n13278 );
    or g4840 ( n8224 , n21924 , n29004 );
    nor g4841 ( n9382 , n25228 , n2160 );
    or g4842 ( n8099 , n10320 , n21607 );
    and g4843 ( n21505 , n27003 , n11260 );
    and g4844 ( n1731 , n5602 , n7301 );
    not g4845 ( n9237 , n6401 );
    not g4846 ( n25269 , n3160 );
    not g4847 ( n13207 , n9869 );
    not g4848 ( n27652 , n18744 );
    or g4849 ( n30058 , n21653 , n23731 );
    not g4850 ( n11193 , n30678 );
    not g4851 ( n14286 , n23948 );
    or g4852 ( n28244 , n21195 , n19305 );
    not g4853 ( n30884 , n23649 );
    or g4854 ( n8743 , n10063 , n27140 );
    xnor g4855 ( n26371 , n20780 , n11789 );
    not g4856 ( n8908 , n11782 );
    and g4857 ( n27685 , n16022 , n30855 );
    not g4858 ( n13196 , n16864 );
    not g4859 ( n24640 , n17580 );
    nor g4860 ( n8990 , n26581 , n2767 );
    xnor g4861 ( n22901 , n870 , n4021 );
    or g4862 ( n19197 , n14417 , n1389 );
    not g4863 ( n26399 , n15479 );
    not g4864 ( n8439 , n26233 );
    not g4865 ( n21012 , n10220 );
    not g4866 ( n3879 , n21122 );
    and g4867 ( n29582 , n8276 , n4295 );
    not g4868 ( n12060 , n20397 );
    not g4869 ( n12853 , n18557 );
    not g4870 ( n5712 , n6599 );
    nor g4871 ( n1734 , n27711 , n31314 );
    or g4872 ( n30136 , n9180 , n31151 );
    or g4873 ( n22258 , n10487 , n9986 );
    xnor g4874 ( n6431 , n2725 , n1308 );
    or g4875 ( n18040 , n9424 , n13640 );
    not g4876 ( n11577 , n29591 );
    and g4877 ( n24957 , n6750 , n29774 );
    buf g4878 ( n20233 , n13657 );
    or g4879 ( n12103 , n28095 , n19449 );
    or g4880 ( n5096 , n26993 , n30256 );
    not g4881 ( n30335 , n14144 );
    xnor g4882 ( n17691 , n2924 , n21064 );
    not g4883 ( n8144 , n154 );
    or g4884 ( n10345 , n19210 , n31703 );
    nor g4885 ( n18928 , n24980 , n6664 );
    not g4886 ( n23438 , n1879 );
    xor g4887 ( n4179 , n18233 , n27177 );
    not g4888 ( n25012 , n4949 );
    xnor g4889 ( n16786 , n9375 , n15438 );
    or g4890 ( n22899 , n18463 , n21823 );
    not g4891 ( n21465 , n16059 );
    or g4892 ( n12939 , n18280 , n15627 );
    xnor g4893 ( n3251 , n13917 , n6206 );
    xnor g4894 ( n18682 , n7241 , n17798 );
    not g4895 ( n12200 , n28809 );
    or g4896 ( n26907 , n23777 , n30958 );
    xnor g4897 ( n6535 , n21338 , n31150 );
    xnor g4898 ( n7235 , n29929 , n20799 );
    nor g4899 ( n4348 , n12760 , n17218 );
    and g4900 ( n24340 , n13208 , n12545 );
    and g4901 ( n7374 , n44 , n9564 );
    not g4902 ( n590 , n27885 );
    xnor g4903 ( n23778 , n23306 , n9935 );
    nor g4904 ( n19940 , n4125 , n5077 );
    xnor g4905 ( n3124 , n29758 , n30713 );
    not g4906 ( n17026 , n24773 );
    buf g4907 ( n29542 , n9217 );
    xnor g4908 ( n14252 , n1189 , n19337 );
    and g4909 ( n1106 , n8923 , n5151 );
    not g4910 ( n18483 , n5719 );
    xnor g4911 ( n2711 , n6351 , n2277 );
    xnor g4912 ( n10714 , n26756 , n3070 );
    and g4913 ( n2025 , n14092 , n25642 );
    not g4914 ( n10997 , n10090 );
    and g4915 ( n30959 , n8442 , n5269 );
    and g4916 ( n27627 , n31595 , n15833 );
    not g4917 ( n15331 , n22119 );
    xnor g4918 ( n30448 , n30002 , n3106 );
    or g4919 ( n11365 , n21571 , n6913 );
    not g4920 ( n18655 , n23871 );
    or g4921 ( n15543 , n2206 , n5097 );
    or g4922 ( n11437 , n7728 , n16633 );
    and g4923 ( n8817 , n19022 , n24453 );
    nor g4924 ( n13169 , n7692 , n4750 );
    xnor g4925 ( n31194 , n638 , n13705 );
    or g4926 ( n23662 , n24816 , n27312 );
    not g4927 ( n31080 , n25510 );
    xnor g4928 ( n24558 , n25383 , n11648 );
    xnor g4929 ( n26615 , n31455 , n12318 );
    or g4930 ( n6241 , n22685 , n13282 );
    or g4931 ( n13168 , n11609 , n3988 );
    not g4932 ( n21909 , n15030 );
    and g4933 ( n12294 , n24364 , n20297 );
    and g4934 ( n22291 , n21727 , n1603 );
    xnor g4935 ( n6893 , n7167 , n27104 );
    not g4936 ( n25763 , n10001 );
    and g4937 ( n5808 , n27616 , n27347 );
    xor g4938 ( n20349 , n25003 , n26075 );
    or g4939 ( n28060 , n508 , n4425 );
    and g4940 ( n27072 , n9202 , n26109 );
    and g4941 ( n28758 , n4651 , n13138 );
    and g4942 ( n27662 , n29983 , n6857 );
    or g4943 ( n23405 , n28425 , n17982 );
    xnor g4944 ( n28618 , n9835 , n24137 );
    not g4945 ( n14338 , n16946 );
    and g4946 ( n31931 , n13816 , n28826 );
    not g4947 ( n11867 , n19956 );
    xnor g4948 ( n20740 , n20219 , n29364 );
    not g4949 ( n1798 , n19189 );
    not g4950 ( n19152 , n15343 );
    or g4951 ( n22604 , n15686 , n16931 );
    or g4952 ( n31225 , n12113 , n28062 );
    xnor g4953 ( n9481 , n26322 , n1195 );
    not g4954 ( n25794 , n13354 );
    and g4955 ( n10767 , n12949 , n26978 );
    or g4956 ( n7691 , n22742 , n31613 );
    not g4957 ( n2596 , n21733 );
    not g4958 ( n26591 , n9613 );
    not g4959 ( n21345 , n29764 );
    nor g4960 ( n524 , n3012 , n11617 );
    xnor g4961 ( n21574 , n705 , n24493 );
    nor g4962 ( n31518 , n12566 , n891 );
    not g4963 ( n30517 , n1665 );
    or g4964 ( n21289 , n11866 , n25464 );
    xnor g4965 ( n3255 , n6438 , n23096 );
    and g4966 ( n6746 , n4853 , n13085 );
    not g4967 ( n26706 , n22447 );
    xnor g4968 ( n24222 , n9085 , n28347 );
    not g4969 ( n20565 , n31204 );
    or g4970 ( n20566 , n28227 , n12899 );
    xnor g4971 ( n12768 , n5487 , n31743 );
    and g4972 ( n8630 , n2796 , n24317 );
    or g4973 ( n5404 , n13752 , n1573 );
    or g4974 ( n31576 , n31995 , n31628 );
    not g4975 ( n27782 , n13839 );
    and g4976 ( n11144 , n3813 , n9603 );
    not g4977 ( n4560 , n13566 );
    and g4978 ( n13187 , n20848 , n22244 );
    xnor g4979 ( n17586 , n22317 , n4493 );
    and g4980 ( n22313 , n14051 , n22847 );
    or g4981 ( n14200 , n3559 , n9243 );
    not g4982 ( n30956 , n20218 );
    or g4983 ( n20780 , n31676 , n17532 );
    xnor g4984 ( n10709 , n27065 , n23934 );
    xnor g4985 ( n2933 , n1028 , n27063 );
    not g4986 ( n22881 , n30702 );
    and g4987 ( n12168 , n18045 , n21493 );
    and g4988 ( n18348 , n15868 , n14285 );
    or g4989 ( n25494 , n90 , n63 );
    not g4990 ( n20973 , n10236 );
    xnor g4991 ( n2680 , n6328 , n9380 );
    not g4992 ( n26038 , n4531 );
    xnor g4993 ( n859 , n14229 , n3023 );
    or g4994 ( n1928 , n3286 , n18250 );
    and g4995 ( n14245 , n4302 , n10659 );
    not g4996 ( n2217 , n8698 );
    and g4997 ( n17674 , n18561 , n27873 );
    not g4998 ( n20503 , n17357 );
    not g4999 ( n26162 , n1344 );
    not g5000 ( n20345 , n18502 );
    xnor g5001 ( n16948 , n7764 , n17166 );
    not g5002 ( n18068 , n31111 );
    not g5003 ( n29420 , n23557 );
    not g5004 ( n3240 , n31785 );
    or g5005 ( n8942 , n5056 , n3766 );
    xnor g5006 ( n3186 , n7452 , n3289 );
    and g5007 ( n25036 , n22032 , n22698 );
    nor g5008 ( n1407 , n16181 , n19228 );
    xnor g5009 ( n19273 , n26894 , n17843 );
    not g5010 ( n8960 , n13868 );
    not g5011 ( n1448 , n24131 );
    xnor g5012 ( n2642 , n11980 , n26233 );
    xnor g5013 ( n25469 , n25570 , n11859 );
    xnor g5014 ( n10362 , n11647 , n21694 );
    nor g5015 ( n22744 , n7302 , n9006 );
    or g5016 ( n21348 , n8026 , n25304 );
    xnor g5017 ( n10693 , n11298 , n15130 );
    not g5018 ( n13908 , n12540 );
    xnor g5019 ( n27181 , n23678 , n24056 );
    not g5020 ( n29080 , n26873 );
    or g5021 ( n284 , n25505 , n15393 );
    xnor g5022 ( n30923 , n21676 , n19441 );
    or g5023 ( n26864 , n6608 , n26808 );
    and g5024 ( n2434 , n18206 , n9238 );
    xnor g5025 ( n9689 , n18937 , n21682 );
    or g5026 ( n28647 , n14248 , n15771 );
    xor g5027 ( n2803 , n18438 , n5077 );
    not g5028 ( n14449 , n14155 );
    and g5029 ( n28292 , n227 , n1719 );
    and g5030 ( n3954 , n9694 , n19992 );
    xnor g5031 ( n11131 , n26386 , n15852 );
    and g5032 ( n18308 , n31950 , n14781 );
    xnor g5033 ( n357 , n7819 , n13400 );
    or g5034 ( n19850 , n15556 , n15752 );
    xnor g5035 ( n449 , n26499 , n4266 );
    and g5036 ( n9771 , n13761 , n15356 );
    and g5037 ( n17087 , n11842 , n26802 );
    nor g5038 ( n29521 , n26598 , n15930 );
    xnor g5039 ( n6144 , n17104 , n7705 );
    and g5040 ( n17973 , n25771 , n1358 );
    xnor g5041 ( n29448 , n4194 , n19295 );
    xnor g5042 ( n5183 , n12427 , n19615 );
    or g5043 ( n1256 , n16815 , n13046 );
    not g5044 ( n27162 , n5060 );
    xnor g5045 ( n14707 , n11133 , n20021 );
    or g5046 ( n18222 , n19008 , n27009 );
    xnor g5047 ( n4285 , n31033 , n14816 );
    not g5048 ( n5951 , n19625 );
    or g5049 ( n25022 , n30408 , n557 );
    or g5050 ( n23085 , n7171 , n18313 );
    xnor g5051 ( n11814 , n26702 , n18541 );
    not g5052 ( n21572 , n5996 );
    and g5053 ( n25474 , n9724 , n24600 );
    or g5054 ( n21126 , n7571 , n12114 );
    not g5055 ( n4111 , n9734 );
    or g5056 ( n9896 , n3631 , n26977 );
    or g5057 ( n6857 , n15073 , n20146 );
    or g5058 ( n30059 , n16193 , n12096 );
    not g5059 ( n5720 , n7140 );
    not g5060 ( n16997 , n17941 );
    and g5061 ( n15812 , n22031 , n1195 );
    not g5062 ( n21393 , n4567 );
    xnor g5063 ( n13333 , n15810 , n22104 );
    or g5064 ( n4044 , n28684 , n16396 );
    xnor g5065 ( n22803 , n24845 , n3340 );
    or g5066 ( n6351 , n5383 , n28195 );
    xnor g5067 ( n25337 , n24807 , n31896 );
    or g5068 ( n693 , n4496 , n9719 );
    or g5069 ( n3209 , n25334 , n3428 );
    or g5070 ( n3931 , n14947 , n26129 );
    not g5071 ( n16792 , n1695 );
    nor g5072 ( n25262 , n3912 , n25076 );
    xnor g5073 ( n4235 , n6126 , n24350 );
    not g5074 ( n30744 , n20799 );
    or g5075 ( n3222 , n24838 , n20348 );
    nor g5076 ( n8026 , n21671 , n466 );
    or g5077 ( n12120 , n2785 , n13315 );
    and g5078 ( n230 , n15303 , n6309 );
    xnor g5079 ( n12437 , n23525 , n784 );
    or g5080 ( n1542 , n4410 , n27672 );
    or g5081 ( n18666 , n29173 , n31582 );
    xnor g5082 ( n14718 , n18980 , n205 );
    not g5083 ( n23921 , n29391 );
    or g5084 ( n10338 , n28655 , n17903 );
    not g5085 ( n10876 , n11643 );
    xnor g5086 ( n12462 , n25344 , n11851 );
    not g5087 ( n28930 , n19783 );
    not g5088 ( n21760 , n30862 );
    nor g5089 ( n22517 , n22610 , n16122 );
    not g5090 ( n20981 , n4298 );
    not g5091 ( n19068 , n27390 );
    not g5092 ( n19224 , n31921 );
    or g5093 ( n3253 , n2272 , n31307 );
    or g5094 ( n19053 , n1273 , n11497 );
    xnor g5095 ( n12991 , n2385 , n15547 );
    not g5096 ( n21120 , n17271 );
    and g5097 ( n11919 , n2867 , n25420 );
    xnor g5098 ( n12831 , n3709 , n24289 );
    not g5099 ( n20488 , n11424 );
    or g5100 ( n29271 , n4355 , n11263 );
    buf g5101 ( n26763 , n24431 );
    xnor g5102 ( n25586 , n24009 , n13394 );
    not g5103 ( n5822 , n11771 );
    xnor g5104 ( n22200 , n30849 , n30257 );
    and g5105 ( n25698 , n29415 , n15309 );
    or g5106 ( n9085 , n24368 , n22071 );
    not g5107 ( n1397 , n31968 );
    or g5108 ( n7790 , n26142 , n13031 );
    xnor g5109 ( n25857 , n19029 , n10420 );
    or g5110 ( n11199 , n31993 , n26493 );
    not g5111 ( n9884 , n17582 );
    or g5112 ( n25142 , n29249 , n8120 );
    not g5113 ( n19102 , n8207 );
    and g5114 ( n6360 , n274 , n8963 );
    xnor g5115 ( n11801 , n27314 , n6396 );
    xnor g5116 ( n1065 , n7185 , n24452 );
    xnor g5117 ( n30266 , n3325 , n17805 );
    or g5118 ( n25411 , n3639 , n31260 );
    and g5119 ( n17347 , n9653 , n9424 );
    or g5120 ( n11053 , n16582 , n19009 );
    nor g5121 ( n13416 , n10416 , n7248 );
    not g5122 ( n4942 , n26534 );
    xnor g5123 ( n23319 , n27782 , n18161 );
    not g5124 ( n9079 , n25187 );
    nor g5125 ( n17723 , n22393 , n2535 );
    not g5126 ( n1543 , n22936 );
    nor g5127 ( n30399 , n22248 , n30106 );
    xnor g5128 ( n10880 , n24043 , n28702 );
    and g5129 ( n20638 , n7403 , n3337 );
    or g5130 ( n9385 , n26380 , n30912 );
    xnor g5131 ( n4607 , n22987 , n12092 );
    not g5132 ( n27986 , n24650 );
    or g5133 ( n14621 , n6508 , n1782 );
    not g5134 ( n16685 , n20380 );
    xnor g5135 ( n27070 , n14717 , n8387 );
    and g5136 ( n7091 , n22349 , n13690 );
    or g5137 ( n1930 , n9063 , n14367 );
    and g5138 ( n11902 , n15108 , n17368 );
    not g5139 ( n2781 , n17110 );
    not g5140 ( n18241 , n15109 );
    or g5141 ( n10162 , n3811 , n6877 );
    not g5142 ( n794 , n4854 );
    or g5143 ( n31556 , n8177 , n26144 );
    or g5144 ( n2946 , n29443 , n26930 );
    and g5145 ( n62 , n22644 , n21269 );
    and g5146 ( n5106 , n4162 , n5553 );
    and g5147 ( n29342 , n19171 , n27525 );
    not g5148 ( n18103 , n22077 );
    not g5149 ( n19298 , n11355 );
    not g5150 ( n23862 , n6766 );
    and g5151 ( n16367 , n15543 , n31594 );
    and g5152 ( n29362 , n8533 , n3468 );
    not g5153 ( n11537 , n18871 );
    or g5154 ( n15814 , n9426 , n20152 );
    and g5155 ( n9372 , n16313 , n10676 );
    and g5156 ( n6573 , n17583 , n26516 );
    not g5157 ( n1098 , n23707 );
    xnor g5158 ( n15048 , n30425 , n17109 );
    or g5159 ( n23656 , n25320 , n28269 );
    xnor g5160 ( n25513 , n18391 , n31773 );
    xnor g5161 ( n12497 , n30326 , n29153 );
    xnor g5162 ( n9572 , n28129 , n27721 );
    not g5163 ( n7813 , n19400 );
    or g5164 ( n7320 , n11278 , n25128 );
    or g5165 ( n250 , n3716 , n14252 );
    and g5166 ( n8286 , n10655 , n28875 );
    not g5167 ( n29825 , n24439 );
    not g5168 ( n15113 , n28827 );
    or g5169 ( n16585 , n28091 , n11958 );
    or g5170 ( n5207 , n28434 , n17179 );
    not g5171 ( n1986 , n9318 );
    nor g5172 ( n13901 , n21520 , n29028 );
    xnor g5173 ( n29520 , n23106 , n16426 );
    not g5174 ( n19172 , n22598 );
    or g5175 ( n27707 , n11201 , n25593 );
    not g5176 ( n28351 , n1665 );
    or g5177 ( n25776 , n138 , n18391 );
    or g5178 ( n17296 , n163 , n31979 );
    not g5179 ( n2522 , n30526 );
    not g5180 ( n26628 , n19615 );
    xnor g5181 ( n16656 , n30325 , n7285 );
    not g5182 ( n23646 , n23112 );
    not g5183 ( n7534 , n30622 );
    or g5184 ( n11384 , n26114 , n2872 );
    xnor g5185 ( n7553 , n25168 , n10305 );
    not g5186 ( n27332 , n13642 );
    and g5187 ( n21497 , n28759 , n22572 );
    not g5188 ( n18439 , n21252 );
    xnor g5189 ( n14527 , n10337 , n30719 );
    not g5190 ( n2027 , n7290 );
    xnor g5191 ( n3460 , n20829 , n7779 );
    not g5192 ( n28426 , n31975 );
    not g5193 ( n26315 , n18557 );
    not g5194 ( n3664 , n18512 );
    or g5195 ( n6740 , n24407 , n23022 );
    or g5196 ( n9665 , n20878 , n26668 );
    nor g5197 ( n4447 , n12600 , n4421 );
    and g5198 ( n28465 , n13070 , n585 );
    or g5199 ( n8589 , n24921 , n15088 );
    and g5200 ( n5694 , n11602 , n31844 );
    or g5201 ( n9573 , n256 , n25016 );
    or g5202 ( n19787 , n13449 , n866 );
    and g5203 ( n12149 , n2425 , n9553 );
    not g5204 ( n21280 , n27501 );
    xnor g5205 ( n22093 , n30145 , n31957 );
    or g5206 ( n25256 , n11182 , n27388 );
    xnor g5207 ( n24180 , n9514 , n10429 );
    xnor g5208 ( n2405 , n4044 , n20570 );
    not g5209 ( n21914 , n5838 );
    nor g5210 ( n16185 , n3508 , n21654 );
    not g5211 ( n14005 , n22664 );
    and g5212 ( n20126 , n21747 , n27114 );
    xnor g5213 ( n6824 , n12731 , n28386 );
    and g5214 ( n17794 , n30927 , n19211 );
    nor g5215 ( n10887 , n10985 , n12773 );
    or g5216 ( n6443 , n6297 , n1641 );
    or g5217 ( n22722 , n8302 , n25114 );
    and g5218 ( n14740 , n8634 , n22495 );
    xnor g5219 ( n10115 , n24865 , n6386 );
    and g5220 ( n19319 , n12258 , n17588 );
    and g5221 ( n8970 , n6538 , n15522 );
    nor g5222 ( n26909 , n21963 , n13496 );
    or g5223 ( n24619 , n13917 , n26484 );
    or g5224 ( n13586 , n13524 , n3581 );
    not g5225 ( n6034 , n12627 );
    xnor g5226 ( n6401 , n15218 , n14308 );
    nor g5227 ( n13793 , n4747 , n2095 );
    xnor g5228 ( n10306 , n29329 , n28047 );
    not g5229 ( n10027 , n12774 );
    xnor g5230 ( n7202 , n7843 , n30227 );
    xnor g5231 ( n10775 , n7705 , n13454 );
    xnor g5232 ( n4342 , n18898 , n14591 );
    not g5233 ( n24288 , n11363 );
    or g5234 ( n28722 , n26456 , n12514 );
    xnor g5235 ( n12380 , n29043 , n8666 );
    and g5236 ( n19778 , n22694 , n17301 );
    or g5237 ( n27406 , n27460 , n7618 );
    or g5238 ( n22273 , n25574 , n11625 );
    and g5239 ( n3684 , n29752 , n24759 );
    not g5240 ( n24409 , n26072 );
    and g5241 ( n30547 , n23214 , n2441 );
    or g5242 ( n21936 , n4153 , n3889 );
    not g5243 ( n9016 , n23562 );
    or g5244 ( n19164 , n818 , n18092 );
    xnor g5245 ( n11056 , n23698 , n18010 );
    and g5246 ( n15402 , n8551 , n31660 );
    and g5247 ( n19269 , n13038 , n12566 );
    or g5248 ( n25850 , n13528 , n5102 );
    not g5249 ( n3912 , n7200 );
    or g5250 ( n10972 , n14612 , n26399 );
    not g5251 ( n5086 , n13930 );
    or g5252 ( n14849 , n4776 , n980 );
    nor g5253 ( n22887 , n451 , n2183 );
    and g5254 ( n24625 , n29627 , n2472 );
    not g5255 ( n25554 , n29259 );
    and g5256 ( n3846 , n21714 , n31072 );
    not g5257 ( n14542 , n5428 );
    and g5258 ( n16650 , n30514 , n15588 );
    or g5259 ( n9631 , n5954 , n28017 );
    not g5260 ( n29259 , n27139 );
    not g5261 ( n16291 , n20403 );
    xor g5262 ( n842 , n28108 , n25195 );
    xnor g5263 ( n22763 , n16248 , n757 );
    and g5264 ( n28080 , n29402 , n13629 );
    and g5265 ( n20824 , n22391 , n25811 );
    not g5266 ( n14516 , n4928 );
    not g5267 ( n17620 , n3408 );
    and g5268 ( n29776 , n31692 , n1747 );
    buf g5269 ( n26006 , n474 );
    xnor g5270 ( n6440 , n28196 , n25519 );
    nor g5271 ( n13979 , n2924 , n8166 );
    or g5272 ( n13217 , n15237 , n5651 );
    not g5273 ( n18237 , n19044 );
    not g5274 ( n27531 , n5794 );
    or g5275 ( n13460 , n7765 , n16720 );
    xnor g5276 ( n26492 , n13194 , n25974 );
    or g5277 ( n19691 , n21083 , n195 );
    buf g5278 ( n22244 , n21246 );
    xnor g5279 ( n30359 , n11462 , n3432 );
    xnor g5280 ( n7444 , n18482 , n20669 );
    xnor g5281 ( n3426 , n26058 , n23739 );
    not g5282 ( n5992 , n9172 );
    not g5283 ( n31921 , n8424 );
    and g5284 ( n22077 , n18324 , n7936 );
    or g5285 ( n13100 , n6352 , n8299 );
    buf g5286 ( n15266 , n5753 );
    and g5287 ( n18860 , n24683 , n5832 );
    or g5288 ( n8070 , n31521 , n10449 );
    not g5289 ( n6667 , n8333 );
    or g5290 ( n1509 , n2278 , n1108 );
    not g5291 ( n15776 , n5069 );
    and g5292 ( n21644 , n5132 , n22045 );
    and g5293 ( n5178 , n13198 , n13176 );
    and g5294 ( n14224 , n23436 , n9470 );
    and g5295 ( n6187 , n12218 , n25839 );
    xnor g5296 ( n25755 , n12551 , n5349 );
    and g5297 ( n2102 , n15244 , n7202 );
    or g5298 ( n2745 , n4019 , n13303 );
    and g5299 ( n11528 , n31273 , n1149 );
    xnor g5300 ( n8326 , n1758 , n14560 );
    xnor g5301 ( n3814 , n6854 , n13270 );
    not g5302 ( n18076 , n25991 );
    not g5303 ( n18610 , n23260 );
    nor g5304 ( n19735 , n9336 , n22977 );
    not g5305 ( n17755 , n14345 );
    not g5306 ( n21818 , n6197 );
    and g5307 ( n9304 , n16375 , n7280 );
    or g5308 ( n23972 , n16600 , n28442 );
    not g5309 ( n9914 , n28438 );
    not g5310 ( n12138 , n8641 );
    xnor g5311 ( n28646 , n30780 , n10445 );
    or g5312 ( n13015 , n4260 , n9060 );
    or g5313 ( n24438 , n950 , n31454 );
    nor g5314 ( n19079 , n11658 , n7314 );
    or g5315 ( n30107 , n31261 , n31745 );
    xor g5316 ( n10067 , n29570 , n20736 );
    nor g5317 ( n772 , n8450 , n1872 );
    and g5318 ( n2379 , n22479 , n7989 );
    or g5319 ( n11134 , n23145 , n13250 );
    not g5320 ( n14411 , n7662 );
    not g5321 ( n31898 , n3313 );
    xnor g5322 ( n19256 , n29874 , n1335 );
    and g5323 ( n15654 , n17273 , n5776 );
    and g5324 ( n15386 , n13182 , n15908 );
    not g5325 ( n4322 , n14876 );
    or g5326 ( n26249 , n28983 , n11466 );
    and g5327 ( n26709 , n29 , n27011 );
    or g5328 ( n27338 , n936 , n27722 );
    xnor g5329 ( n29457 , n20155 , n11373 );
    xnor g5330 ( n28347 , n26331 , n9751 );
    not g5331 ( n13501 , n1241 );
    not g5332 ( n10504 , n30908 );
    or g5333 ( n6156 , n4208 , n30933 );
    xnor g5334 ( n1636 , n24512 , n10474 );
    xnor g5335 ( n30164 , n20905 , n22434 );
    not g5336 ( n16115 , n28720 );
    xnor g5337 ( n684 , n10436 , n19706 );
    and g5338 ( n7827 , n20130 , n24350 );
    or g5339 ( n24780 , n21888 , n268 );
    xnor g5340 ( n159 , n2369 , n25580 );
    and g5341 ( n15816 , n23179 , n15749 );
    and g5342 ( n23261 , n26293 , n17935 );
    or g5343 ( n10448 , n28557 , n31912 );
    nor g5344 ( n1540 , n6349 , n30189 );
    nor g5345 ( n20907 , n24907 , n21488 );
    xnor g5346 ( n10498 , n8220 , n3131 );
    or g5347 ( n6765 , n4047 , n23488 );
    xnor g5348 ( n30567 , n24484 , n764 );
    xnor g5349 ( n18812 , n21532 , n7771 );
    nor g5350 ( n8020 , n3987 , n24273 );
    and g5351 ( n28761 , n16486 , n8294 );
    xnor g5352 ( n3731 , n15953 , n10677 );
    or g5353 ( n29532 , n20038 , n26207 );
    or g5354 ( n10582 , n30457 , n16182 );
    not g5355 ( n23966 , n23344 );
    not g5356 ( n14694 , n15829 );
    and g5357 ( n24318 , n23325 , n28556 );
    xor g5358 ( n13083 , n30292 , n25758 );
    and g5359 ( n21704 , n21220 , n4897 );
    not g5360 ( n10938 , n3618 );
    or g5361 ( n7073 , n17168 , n12579 );
    nor g5362 ( n10908 , n18490 , n10967 );
    not g5363 ( n27930 , n20175 );
    and g5364 ( n15652 , n23995 , n20881 );
    xnor g5365 ( n28583 , n5079 , n17325 );
    or g5366 ( n4646 , n13535 , n26753 );
    xnor g5367 ( n776 , n28006 , n508 );
    xnor g5368 ( n16225 , n2180 , n17557 );
    or g5369 ( n12021 , n23601 , n11022 );
    not g5370 ( n16364 , n31672 );
    or g5371 ( n5931 , n12252 , n29479 );
    not g5372 ( n9987 , n14489 );
    or g5373 ( n17465 , n1267 , n29607 );
    not g5374 ( n20344 , n7262 );
    or g5375 ( n7072 , n2525 , n27991 );
    not g5376 ( n18821 , n15756 );
    not g5377 ( n31283 , n21781 );
    xnor g5378 ( n22913 , n7555 , n11761 );
    nor g5379 ( n19032 , n21185 , n27805 );
    buf g5380 ( n22349 , n16448 );
    and g5381 ( n15000 , n23111 , n23127 );
    or g5382 ( n9780 , n30185 , n31538 );
    or g5383 ( n17889 , n25315 , n19664 );
    not g5384 ( n7004 , n15639 );
    xnor g5385 ( n10405 , n12331 , n29604 );
    xnor g5386 ( n17760 , n8878 , n17755 );
    not g5387 ( n1384 , n4924 );
    not g5388 ( n21248 , n18598 );
    nor g5389 ( n15860 , n11738 , n26185 );
    not g5390 ( n13017 , n16697 );
    xnor g5391 ( n18449 , n26864 , n9449 );
    not g5392 ( n8110 , n31973 );
    and g5393 ( n17807 , n4882 , n209 );
    xnor g5394 ( n1906 , n15616 , n1147 );
    not g5395 ( n20790 , n11711 );
    xnor g5396 ( n2358 , n3972 , n18298 );
    not g5397 ( n15672 , n21033 );
    xnor g5398 ( n31927 , n13431 , n28063 );
    xnor g5399 ( n25189 , n18574 , n25125 );
    or g5400 ( n8307 , n24228 , n20470 );
    xnor g5401 ( n24322 , n29221 , n888 );
    xnor g5402 ( n11956 , n8549 , n11574 );
    xnor g5403 ( n20447 , n29335 , n2150 );
    not g5404 ( n27020 , n20274 );
    or g5405 ( n7536 , n24226 , n7068 );
    xnor g5406 ( n18633 , n19991 , n30360 );
    nor g5407 ( n20104 , n4220 , n27855 );
    xnor g5408 ( n3829 , n18436 , n17060 );
    xnor g5409 ( n27179 , n16092 , n27064 );
    xnor g5410 ( n24909 , n11939 , n1708 );
    or g5411 ( n6817 , n30658 , n24876 );
    not g5412 ( n6053 , n18442 );
    nor g5413 ( n1421 , n24512 , n2813 );
    not g5414 ( n7379 , n7593 );
    or g5415 ( n29973 , n13166 , n29103 );
    and g5416 ( n13804 , n13880 , n12819 );
    buf g5417 ( n21464 , n19642 );
    not g5418 ( n19478 , n25819 );
    xnor g5419 ( n18022 , n21029 , n26732 );
    not g5420 ( n5500 , n14375 );
    not g5421 ( n15623 , n17979 );
    or g5422 ( n13427 , n25452 , n29172 );
    and g5423 ( n29791 , n13390 , n31223 );
    nor g5424 ( n31862 , n9116 , n25810 );
    xnor g5425 ( n5723 , n13312 , n14450 );
    not g5426 ( n23855 , n14556 );
    not g5427 ( n15373 , n28273 );
    not g5428 ( n24732 , n19314 );
    xnor g5429 ( n14171 , n30900 , n22141 );
    xnor g5430 ( n7540 , n9747 , n31440 );
    or g5431 ( n25249 , n20850 , n1711 );
    or g5432 ( n3704 , n20095 , n4486 );
    and g5433 ( n29828 , n21481 , n21738 );
    not g5434 ( n20150 , n28781 );
    nor g5435 ( n12023 , n15997 , n3014 );
    or g5436 ( n4991 , n27554 , n29671 );
    or g5437 ( n12818 , n10490 , n6416 );
    nor g5438 ( n20944 , n5628 , n18913 );
    nor g5439 ( n5359 , n21603 , n9312 );
    and g5440 ( n10652 , n12051 , n31664 );
    not g5441 ( n12898 , n11462 );
    not g5442 ( n11202 , n26751 );
    and g5443 ( n8470 , n30352 , n30792 );
    not g5444 ( n14498 , n21302 );
    not g5445 ( n28597 , n22533 );
    xnor g5446 ( n25519 , n5567 , n13634 );
    or g5447 ( n7633 , n16219 , n30166 );
    or g5448 ( n11652 , n6425 , n1623 );
    not g5449 ( n13170 , n6938 );
    and g5450 ( n22537 , n26501 , n20530 );
    or g5451 ( n17936 , n2895 , n13713 );
    buf g5452 ( n22345 , n8253 );
    nor g5453 ( n2966 , n14795 , n22866 );
    not g5454 ( n4617 , n5380 );
    or g5455 ( n6318 , n5289 , n31804 );
    not g5456 ( n27710 , n986 );
    or g5457 ( n9128 , n15009 , n18921 );
    not g5458 ( n6553 , n27971 );
    not g5459 ( n25260 , n22418 );
    xnor g5460 ( n24147 , n22204 , n3157 );
    not g5461 ( n14249 , n5654 );
    or g5462 ( n11282 , n17628 , n11801 );
    or g5463 ( n27616 , n30874 , n30304 );
    or g5464 ( n15175 , n17185 , n22536 );
    xor g5465 ( n401 , n4837 , n5458 );
    or g5466 ( n19650 , n26171 , n3052 );
    nor g5467 ( n16528 , n12433 , n4229 );
    and g5468 ( n16820 , n28530 , n25034 );
    and g5469 ( n15545 , n20112 , n17765 );
    not g5470 ( n12994 , n20877 );
    or g5471 ( n21037 , n15 , n26454 );
    nor g5472 ( n4522 , n27501 , n2849 );
    or g5473 ( n20911 , n5529 , n6654 );
    xnor g5474 ( n527 , n11767 , n25068 );
    xnor g5475 ( n1888 , n16658 , n13351 );
    not g5476 ( n11054 , n23415 );
    xnor g5477 ( n6554 , n2657 , n31792 );
    not g5478 ( n5596 , n16075 );
    xnor g5479 ( n24929 , n18291 , n18159 );
    not g5480 ( n19510 , n10635 );
    nor g5481 ( n5689 , n28192 , n11332 );
    and g5482 ( n15912 , n30215 , n24753 );
    buf g5483 ( n22104 , n31575 );
    xnor g5484 ( n3194 , n8739 , n30574 );
    xnor g5485 ( n323 , n24157 , n13785 );
    or g5486 ( n13750 , n6141 , n25864 );
    or g5487 ( n12592 , n17791 , n9668 );
    and g5488 ( n8465 , n20559 , n24915 );
    or g5489 ( n24359 , n23960 , n21019 );
    or g5490 ( n24637 , n3724 , n18333 );
    xor g5491 ( n17042 , n27647 , n28942 );
    and g5492 ( n9101 , n2805 , n19509 );
    not g5493 ( n10769 , n7904 );
    not g5494 ( n15735 , n1318 );
    not g5495 ( n30182 , n28524 );
    xnor g5496 ( n19287 , n31031 , n17284 );
    not g5497 ( n29507 , n4908 );
    nor g5498 ( n347 , n27355 , n19274 );
    and g5499 ( n5092 , n16428 , n10054 );
    and g5500 ( n10856 , n22233 , n31060 );
    xnor g5501 ( n15370 , n8988 , n7046 );
    and g5502 ( n23765 , n18300 , n27643 );
    not g5503 ( n26321 , n7592 );
    nor g5504 ( n5307 , n5948 , n12489 );
    and g5505 ( n9946 , n17474 , n12857 );
    xnor g5506 ( n16714 , n9792 , n15669 );
    nor g5507 ( n4514 , n24969 , n1957 );
    not g5508 ( n21447 , n2558 );
    not g5509 ( n282 , n5290 );
    nor g5510 ( n27125 , n7543 , n28197 );
    nor g5511 ( n3232 , n10088 , n28020 );
    not g5512 ( n1077 , n12036 );
    nor g5513 ( n31959 , n26832 , n21259 );
    not g5514 ( n27244 , n11005 );
    or g5515 ( n3923 , n4793 , n1463 );
    xnor g5516 ( n16187 , n10230 , n4199 );
    xnor g5517 ( n11016 , n29865 , n31579 );
    xnor g5518 ( n9537 , n17532 , n10334 );
    not g5519 ( n26210 , n16791 );
    or g5520 ( n26727 , n8351 , n2774 );
    xnor g5521 ( n31344 , n14743 , n667 );
    and g5522 ( n15299 , n7334 , n30512 );
    or g5523 ( n17698 , n22139 , n18240 );
    not g5524 ( n8075 , n16478 );
    xnor g5525 ( n13230 , n11362 , n8989 );
    not g5526 ( n23731 , n8939 );
    not g5527 ( n25929 , n15 );
    and g5528 ( n19672 , n20689 , n19053 );
    and g5529 ( n12557 , n23520 , n1025 );
    not g5530 ( n4601 , n27327 );
    not g5531 ( n22640 , n2937 );
    or g5532 ( n28561 , n11688 , n9284 );
    or g5533 ( n8772 , n2394 , n18560 );
    and g5534 ( n17268 , n23140 , n22999 );
    xnor g5535 ( n3786 , n16906 , n3405 );
    and g5536 ( n29094 , n2902 , n24278 );
    xnor g5537 ( n11264 , n18158 , n5168 );
    xnor g5538 ( n19435 , n4350 , n24056 );
    not g5539 ( n26220 , n15261 );
    xnor g5540 ( n26633 , n6892 , n6931 );
    or g5541 ( n15443 , n6055 , n12904 );
    not g5542 ( n10053 , n31043 );
    nor g5543 ( n9902 , n11309 , n3959 );
    or g5544 ( n17643 , n7350 , n4338 );
    xor g5545 ( n27917 , n17549 , n16201 );
    and g5546 ( n17326 , n22946 , n2085 );
    xnor g5547 ( n24786 , n22193 , n3820 );
    xnor g5548 ( n15858 , n18281 , n13506 );
    or g5549 ( n13361 , n8565 , n14125 );
    or g5550 ( n19265 , n23361 , n13622 );
    not g5551 ( n1632 , n31470 );
    or g5552 ( n3373 , n1053 , n8127 );
    or g5553 ( n31838 , n25659 , n14295 );
    or g5554 ( n27174 , n1032 , n19093 );
    and g5555 ( n27402 , n4259 , n26307 );
    not g5556 ( n3212 , n6797 );
    not g5557 ( n18795 , n16298 );
    not g5558 ( n7453 , n7958 );
    nor g5559 ( n22373 , n5113 , n22470 );
    not g5560 ( n12306 , n21408 );
    not g5561 ( n21897 , n7014 );
    and g5562 ( n9621 , n9584 , n2396 );
    not g5563 ( n8182 , n5664 );
    xnor g5564 ( n20309 , n615 , n9487 );
    or g5565 ( n8777 , n8490 , n22770 );
    xnor g5566 ( n27413 , n23195 , n29569 );
    and g5567 ( n14296 , n22477 , n27977 );
    not g5568 ( n10772 , n10139 );
    xnor g5569 ( n31078 , n14219 , n4847 );
    not g5570 ( n2831 , n17750 );
    not g5571 ( n4539 , n24857 );
    not g5572 ( n2089 , n11321 );
    xnor g5573 ( n10083 , n14304 , n14401 );
    not g5574 ( n14037 , n28112 );
    or g5575 ( n19718 , n1570 , n30115 );
    or g5576 ( n20440 , n15568 , n4750 );
    or g5577 ( n25784 , n22319 , n26029 );
    not g5578 ( n10038 , n2205 );
    not g5579 ( n754 , n20789 );
    not g5580 ( n19561 , n11262 );
    not g5581 ( n19364 , n1293 );
    or g5582 ( n6541 , n31331 , n27484 );
    or g5583 ( n26276 , n19965 , n5604 );
    not g5584 ( n304 , n4700 );
    or g5585 ( n15777 , n18115 , n25955 );
    not g5586 ( n16925 , n23037 );
    nor g5587 ( n26886 , n21963 , n21441 );
    xnor g5588 ( n24652 , n4122 , n25585 );
    or g5589 ( n13608 , n16370 , n23015 );
    buf g5590 ( n22522 , n23757 );
    xnor g5591 ( n5734 , n3122 , n6560 );
    or g5592 ( n14820 , n5621 , n31005 );
    not g5593 ( n31572 , n1234 );
    nor g5594 ( n2189 , n8029 , n3140 );
    and g5595 ( n5529 , n11050 , n664 );
    not g5596 ( n18577 , n20864 );
    nor g5597 ( n10560 , n5241 , n15664 );
    not g5598 ( n2866 , n18449 );
    not g5599 ( n10989 , n8221 );
    xnor g5600 ( n18873 , n9441 , n4536 );
    or g5601 ( n23985 , n17836 , n29719 );
    not g5602 ( n9862 , n20392 );
    or g5603 ( n31136 , n13419 , n27965 );
    nor g5604 ( n12237 , n11361 , n19185 );
    not g5605 ( n23829 , n5392 );
    nor g5606 ( n28673 , n22546 , n15939 );
    nor g5607 ( n26822 , n2001 , n14636 );
    and g5608 ( n28834 , n20702 , n13059 );
    not g5609 ( n6135 , n29550 );
    not g5610 ( n30775 , n28372 );
    xnor g5611 ( n13461 , n16959 , n29589 );
    not g5612 ( n19372 , n5733 );
    and g5613 ( n9031 , n16804 , n27976 );
    xnor g5614 ( n21580 , n22086 , n24416 );
    not g5615 ( n6230 , n30999 );
    not g5616 ( n5503 , n14983 );
    not g5617 ( n23394 , n7345 );
    and g5618 ( n7145 , n1587 , n29993 );
    not g5619 ( n28655 , n23552 );
    or g5620 ( n28848 , n15749 , n26787 );
    or g5621 ( n25619 , n13125 , n2768 );
    or g5622 ( n19018 , n26259 , n798 );
    and g5623 ( n14055 , n22065 , n16078 );
    and g5624 ( n27293 , n6059 , n12843 );
    not g5625 ( n12541 , n31491 );
    nor g5626 ( n21306 , n30505 , n29075 );
    and g5627 ( n23915 , n13950 , n6926 );
    not g5628 ( n29519 , n8808 );
    xnor g5629 ( n16603 , n816 , n31772 );
    or g5630 ( n14051 , n30399 , n13396 );
    xnor g5631 ( n27298 , n9414 , n3307 );
    xnor g5632 ( n10282 , n18312 , n31019 );
    or g5633 ( n16749 , n5307 , n21828 );
    nor g5634 ( n21201 , n17108 , n5082 );
    xnor g5635 ( n4471 , n11648 , n20390 );
    xnor g5636 ( n27313 , n17737 , n28642 );
    xnor g5637 ( n19117 , n2534 , n5998 );
    not g5638 ( n11225 , n20066 );
    xnor g5639 ( n28105 , n22861 , n15924 );
    xnor g5640 ( n26729 , n24529 , n4056 );
    or g5641 ( n11243 , n18551 , n23786 );
    or g5642 ( n24543 , n7096 , n22752 );
    not g5643 ( n5082 , n19117 );
    nor g5644 ( n12180 , n1923 , n17923 );
    xnor g5645 ( n20029 , n1697 , n21097 );
    xnor g5646 ( n10764 , n16831 , n19250 );
    and g5647 ( n5741 , n14626 , n24553 );
    xnor g5648 ( n29393 , n24973 , n17461 );
    nor g5649 ( n4501 , n11984 , n9964 );
    not g5650 ( n26558 , n6354 );
    not g5651 ( n32009 , n29834 );
    not g5652 ( n22974 , n5108 );
    and g5653 ( n30611 , n6264 , n23355 );
    nor g5654 ( n31001 , n825 , n18974 );
    and g5655 ( n23883 , n18563 , n14968 );
    or g5656 ( n5235 , n14690 , n18264 );
    nor g5657 ( n16237 , n8042 , n12001 );
    not g5658 ( n25335 , n1337 );
    xnor g5659 ( n23530 , n22617 , n10403 );
    xnor g5660 ( n14584 , n13606 , n14515 );
    xnor g5661 ( n12243 , n3146 , n29522 );
    xnor g5662 ( n2195 , n5710 , n21708 );
    xnor g5663 ( n4843 , n31359 , n25805 );
    and g5664 ( n15485 , n6047 , n11162 );
    or g5665 ( n24930 , n30357 , n29544 );
    not g5666 ( n5982 , n23463 );
    not g5667 ( n956 , n2883 );
    not g5668 ( n25837 , n9353 );
    xnor g5669 ( n17171 , n14839 , n2200 );
    or g5670 ( n313 , n917 , n20873 );
    or g5671 ( n3150 , n17235 , n17127 );
    nor g5672 ( n3785 , n27235 , n30277 );
    and g5673 ( n24993 , n8202 , n30977 );
    not g5674 ( n24893 , n15999 );
    or g5675 ( n21224 , n26974 , n4511 );
    and g5676 ( n2875 , n18343 , n23975 );
    xnor g5677 ( n22940 , n28413 , n7651 );
    and g5678 ( n25847 , n13827 , n21512 );
    or g5679 ( n4302 , n25639 , n4354 );
    xnor g5680 ( n5510 , n20700 , n16597 );
    not g5681 ( n27733 , n12730 );
    and g5682 ( n9095 , n22560 , n31261 );
    not g5683 ( n15076 , n29315 );
    and g5684 ( n19176 , n14920 , n22762 );
    and g5685 ( n8595 , n27222 , n16405 );
    and g5686 ( n14916 , n3395 , n4214 );
    nor g5687 ( n30278 , n21324 , n9753 );
    not g5688 ( n31982 , n3506 );
    xnor g5689 ( n21124 , n21074 , n10031 );
    and g5690 ( n3092 , n2944 , n24861 );
    buf g5691 ( n13764 , n26130 );
    xnor g5692 ( n28009 , n29352 , n9978 );
    or g5693 ( n29757 , n11169 , n26869 );
    nor g5694 ( n14732 , n18929 , n11168 );
    not g5695 ( n11554 , n26122 );
    xnor g5696 ( n8323 , n22283 , n21580 );
    not g5697 ( n15731 , n5953 );
    xnor g5698 ( n904 , n24152 , n26004 );
    or g5699 ( n12332 , n12806 , n13514 );
    nor g5700 ( n2770 , n29059 , n4009 );
    and g5701 ( n9756 , n23807 , n2094 );
    and g5702 ( n27192 , n25893 , n14036 );
    or g5703 ( n23286 , n19003 , n7092 );
    or g5704 ( n1164 , n2797 , n17662 );
    or g5705 ( n1038 , n25102 , n7835 );
    xor g5706 ( n13808 , n8785 , n19666 );
    not g5707 ( n5350 , n10044 );
    nor g5708 ( n27709 , n3588 , n4287 );
    or g5709 ( n9742 , n6343 , n24888 );
    not g5710 ( n17648 , n20677 );
    or g5711 ( n5601 , n19735 , n7704 );
    not g5712 ( n12065 , n20708 );
    nor g5713 ( n9120 , n7466 , n18743 );
    nor g5714 ( n20776 , n31366 , n15436 );
    xnor g5715 ( n16562 , n6479 , n3843 );
    xnor g5716 ( n25934 , n7804 , n24983 );
    or g5717 ( n5497 , n6696 , n10943 );
    xnor g5718 ( n14066 , n16558 , n10334 );
    or g5719 ( n17411 , n20664 , n22115 );
    not g5720 ( n29120 , n13886 );
    xnor g5721 ( n14271 , n26371 , n9043 );
    and g5722 ( n26170 , n14278 , n21868 );
    or g5723 ( n25888 , n22408 , n29817 );
    or g5724 ( n23745 , n20632 , n22924 );
    xnor g5725 ( n8680 , n2517 , n10705 );
    or g5726 ( n3832 , n18243 , n17547 );
    nor g5727 ( n30322 , n9702 , n31247 );
    not g5728 ( n6679 , n21447 );
    or g5729 ( n24508 , n23703 , n11572 );
    or g5730 ( n19947 , n9136 , n5496 );
    not g5731 ( n8520 , n17667 );
    not g5732 ( n3691 , n24066 );
    not g5733 ( n3792 , n30761 );
    or g5734 ( n22674 , n4257 , n12125 );
    not g5735 ( n11427 , n7230 );
    not g5736 ( n22154 , n469 );
    or g5737 ( n8828 , n31099 , n23877 );
    xor g5738 ( n288 , n91 , n19481 );
    not g5739 ( n28241 , n26082 );
    and g5740 ( n31620 , n5754 , n14848 );
    xnor g5741 ( n11471 , n18025 , n25333 );
    xnor g5742 ( n5662 , n17109 , n7593 );
    nor g5743 ( n15013 , n22615 , n24141 );
    or g5744 ( n10782 , n19675 , n22371 );
    not g5745 ( n11962 , n30898 );
    or g5746 ( n23412 , n9192 , n23781 );
    not g5747 ( n17339 , n11373 );
    and g5748 ( n22046 , n3658 , n25583 );
    not g5749 ( n4173 , n2562 );
    not g5750 ( n26824 , n21574 );
    nor g5751 ( n20147 , n16075 , n17235 );
    xnor g5752 ( n4288 , n312 , n26549 );
    not g5753 ( n4950 , n20709 );
    and g5754 ( n30759 , n9068 , n3729 );
    not g5755 ( n17756 , n23677 );
    xnor g5756 ( n4995 , n11616 , n23681 );
    and g5757 ( n4572 , n5017 , n6471 );
    nor g5758 ( n6368 , n8283 , n4432 );
    or g5759 ( n23 , n3782 , n26787 );
    or g5760 ( n13550 , n25778 , n18912 );
    or g5761 ( n28530 , n593 , n9583 );
    nor g5762 ( n7822 , n14445 , n2952 );
    not g5763 ( n30258 , n24995 );
    or g5764 ( n10342 , n27645 , n844 );
    not g5765 ( n3902 , n30262 );
    nor g5766 ( n140 , n18930 , n3651 );
    not g5767 ( n16811 , n18795 );
    nor g5768 ( n18963 , n22025 , n26362 );
    or g5769 ( n5756 , n17208 , n18482 );
    and g5770 ( n25711 , n13673 , n11418 );
    or g5771 ( n5903 , n1068 , n20303 );
    nor g5772 ( n19156 , n10196 , n21242 );
    or g5773 ( n1603 , n29079 , n10444 );
    xnor g5774 ( n25924 , n17246 , n7009 );
    not g5775 ( n7978 , n28878 );
    xnor g5776 ( n12009 , n210 , n18686 );
    xnor g5777 ( n12871 , n557 , n20169 );
    xnor g5778 ( n24327 , n11501 , n5409 );
    or g5779 ( n2351 , n3427 , n18327 );
    not g5780 ( n11192 , n2255 );
    or g5781 ( n16573 , n862 , n22044 );
    not g5782 ( n20151 , n5067 );
    xnor g5783 ( n14490 , n25901 , n21844 );
    not g5784 ( n14474 , n11354 );
    and g5785 ( n29852 , n24722 , n6718 );
    not g5786 ( n22039 , n15436 );
    not g5787 ( n18029 , n8995 );
    not g5788 ( n22809 , n4459 );
    not g5789 ( n12642 , n6423 );
    or g5790 ( n12106 , n28483 , n15720 );
    and g5791 ( n29353 , n15967 , n27080 );
    or g5792 ( n23515 , n7593 , n24365 );
    not g5793 ( n30872 , n17954 );
    xnor g5794 ( n25198 , n4162 , n30757 );
    and g5795 ( n15996 , n14709 , n17692 );
    and g5796 ( n15070 , n10963 , n20091 );
    and g5797 ( n1907 , n26127 , n31508 );
    xnor g5798 ( n22453 , n4047 , n10847 );
    xnor g5799 ( n15213 , n24264 , n27187 );
    and g5800 ( n25059 , n18288 , n2800 );
    not g5801 ( n6791 , n25242 );
    or g5802 ( n13369 , n2876 , n22721 );
    not g5803 ( n7676 , n6160 );
    nor g5804 ( n11174 , n17515 , n5098 );
    xnor g5805 ( n24286 , n27534 , n10981 );
    or g5806 ( n2481 , n1442 , n14685 );
    not g5807 ( n20322 , n17271 );
    not g5808 ( n26537 , n28185 );
    xnor g5809 ( n17170 , n29952 , n20775 );
    xnor g5810 ( n29406 , n1935 , n24988 );
    not g5811 ( n2813 , n24246 );
    xnor g5812 ( n13981 , n24578 , n20390 );
    nor g5813 ( n7337 , n7696 , n18233 );
    or g5814 ( n31093 , n23130 , n31422 );
    xnor g5815 ( n6409 , n18818 , n24860 );
    not g5816 ( n26225 , n14324 );
    not g5817 ( n15906 , n26294 );
    or g5818 ( n23213 , n6800 , n10835 );
    or g5819 ( n22980 , n3454 , n1687 );
    and g5820 ( n6090 , n28925 , n16245 );
    xnor g5821 ( n18722 , n29282 , n19913 );
    not g5822 ( n18924 , n6698 );
    not g5823 ( n7078 , n1592 );
    xnor g5824 ( n1893 , n30745 , n14754 );
    xnor g5825 ( n26519 , n13732 , n20825 );
    or g5826 ( n22105 , n13188 , n31002 );
    and g5827 ( n24341 , n17203 , n24282 );
    or g5828 ( n160 , n14717 , n26023 );
    or g5829 ( n3851 , n8750 , n3695 );
    not g5830 ( n20058 , n24765 );
    not g5831 ( n9376 , n1132 );
    and g5832 ( n10815 , n3802 , n28990 );
    not g5833 ( n16339 , n11225 );
    or g5834 ( n21555 , n7311 , n27224 );
    xnor g5835 ( n14070 , n27424 , n16030 );
    and g5836 ( n15548 , n23667 , n11065 );
    or g5837 ( n30076 , n20379 , n13580 );
    xnor g5838 ( n28801 , n10718 , n674 );
    or g5839 ( n19104 , n21671 , n31812 );
    and g5840 ( n21367 , n1184 , n20564 );
    not g5841 ( n6171 , n12398 );
    buf g5842 ( n28063 , n6564 );
    xnor g5843 ( n16512 , n25351 , n8114 );
    xnor g5844 ( n6909 , n9318 , n8919 );
    xnor g5845 ( n10623 , n11257 , n2629 );
    xnor g5846 ( n30139 , n25360 , n27805 );
    xnor g5847 ( n24839 , n84 , n6803 );
    nor g5848 ( n14702 , n8713 , n22738 );
    not g5849 ( n20254 , n671 );
    not g5850 ( n10897 , n25689 );
    not g5851 ( n7804 , n25296 );
    nor g5852 ( n15673 , n10624 , n11767 );
    nor g5853 ( n27339 , n14795 , n7316 );
    xnor g5854 ( n21658 , n28557 , n19474 );
    and g5855 ( n13919 , n14748 , n29210 );
    not g5856 ( n25621 , n1945 );
    not g5857 ( n20712 , n11801 );
    not g5858 ( n27853 , n8896 );
    or g5859 ( n10274 , n7791 , n2479 );
    or g5860 ( n11163 , n6978 , n23853 );
    xnor g5861 ( n6666 , n24645 , n16180 );
    or g5862 ( n10597 , n15096 , n6761 );
    xnor g5863 ( n25047 , n9066 , n24712 );
    or g5864 ( n19022 , n5952 , n31423 );
    nor g5865 ( n26149 , n1244 , n6208 );
    nor g5866 ( n25486 , n11132 , n10747 );
    nor g5867 ( n31737 , n21603 , n30936 );
    and g5868 ( n7538 , n8601 , n851 );
    nor g5869 ( n15960 , n8329 , n28007 );
    not g5870 ( n12573 , n9005 );
    and g5871 ( n17192 , n29504 , n25914 );
    or g5872 ( n26071 , n28089 , n5979 );
    xnor g5873 ( n13265 , n27388 , n22509 );
    not g5874 ( n29061 , n18103 );
    not g5875 ( n25187 , n23649 );
    and g5876 ( n13794 , n4635 , n13809 );
    not g5877 ( n19675 , n8713 );
    xnor g5878 ( n15937 , n25029 , n1465 );
    or g5879 ( n28436 , n22146 , n22959 );
    and g5880 ( n6473 , n6994 , n5487 );
    xnor g5881 ( n21664 , n18633 , n31481 );
    buf g5882 ( n16674 , n14835 );
    not g5883 ( n22081 , n29175 );
    not g5884 ( n11048 , n7425 );
    not g5885 ( n29201 , n21793 );
    or g5886 ( n8692 , n30240 , n29408 );
    xnor g5887 ( n19258 , n16099 , n8493 );
    nor g5888 ( n22217 , n4875 , n12263 );
    nor g5889 ( n2560 , n344 , n7641 );
    or g5890 ( n25685 , n20557 , n11156 );
    xnor g5891 ( n23282 , n14904 , n28085 );
    not g5892 ( n8757 , n12812 );
    not g5893 ( n20013 , n6912 );
    xnor g5894 ( n24028 , n24531 , n18829 );
    and g5895 ( n9251 , n14832 , n4357 );
    not g5896 ( n26260 , n2834 );
    xnor g5897 ( n23603 , n9198 , n3234 );
    not g5898 ( n11172 , n16132 );
    not g5899 ( n5498 , n17951 );
    xnor g5900 ( n16420 , n3996 , n9209 );
    and g5901 ( n8101 , n26562 , n1566 );
    or g5902 ( n13679 , n29889 , n18913 );
    not g5903 ( n19198 , n14386 );
    not g5904 ( n25653 , n16411 );
    nor g5905 ( n13798 , n4865 , n3495 );
    or g5906 ( n20596 , n11971 , n6643 );
    not g5907 ( n29319 , n30913 );
    xor g5908 ( n10082 , n16371 , n14703 );
    xnor g5909 ( n16119 , n14363 , n12605 );
    or g5910 ( n22479 , n7711 , n25777 );
    not g5911 ( n18004 , n26237 );
    or g5912 ( n17996 , n30899 , n19812 );
    not g5913 ( n18279 , n17010 );
    nor g5914 ( n15496 , n24086 , n13192 );
    not g5915 ( n6128 , n13509 );
    and g5916 ( n24592 , n23985 , n6023 );
    or g5917 ( n18513 , n7184 , n17837 );
    nor g5918 ( n11991 , n28983 , n10810 );
    not g5919 ( n21277 , n13563 );
    not g5920 ( n11010 , n31822 );
    not g5921 ( n13413 , n2150 );
    or g5922 ( n10968 , n21056 , n30437 );
    not g5923 ( n835 , n21033 );
    not g5924 ( n3636 , n11036 );
    or g5925 ( n12272 , n880 , n20463 );
    not g5926 ( n26349 , n3606 );
    or g5927 ( n13261 , n32007 , n23177 );
    or g5928 ( n15493 , n13741 , n9512 );
    not g5929 ( n9730 , n11070 );
    and g5930 ( n31285 , n9742 , n13015 );
    nor g5931 ( n21218 , n18551 , n15749 );
    nor g5932 ( n11378 , n15436 , n18551 );
    not g5933 ( n8391 , n12571 );
    nor g5934 ( n29373 , n23195 , n13700 );
    or g5935 ( n21635 , n5050 , n2613 );
    nor g5936 ( n27776 , n24964 , n24675 );
    or g5937 ( n13377 , n29782 , n24386 );
    xnor g5938 ( n4005 , n25153 , n4148 );
    nor g5939 ( n1581 , n285 , n23471 );
    or g5940 ( n31040 , n7950 , n15654 );
    not g5941 ( n11566 , n21773 );
    not g5942 ( n1840 , n7890 );
    xnor g5943 ( n4536 , n27962 , n18203 );
    not g5944 ( n13147 , n27186 );
    xnor g5945 ( n31536 , n9448 , n10262 );
    buf g5946 ( n18312 , n19857 );
    nor g5947 ( n23374 , n25343 , n31265 );
    or g5948 ( n17933 , n25504 , n12845 );
    or g5949 ( n11922 , n9181 , n4724 );
    xnor g5950 ( n31979 , n1106 , n17568 );
    nor g5951 ( n6031 , n31722 , n4992 );
    and g5952 ( n28144 , n12405 , n10662 );
    and g5953 ( n22624 , n18737 , n10153 );
    or g5954 ( n5886 , n30128 , n31976 );
    xnor g5955 ( n11627 , n11987 , n13264 );
    not g5956 ( n22734 , n14421 );
    or g5957 ( n8406 , n20024 , n22892 );
    or g5958 ( n6557 , n531 , n26128 );
    and g5959 ( n25867 , n23831 , n11568 );
    not g5960 ( n30663 , n5749 );
    xnor g5961 ( n29084 , n13919 , n19998 );
    or g5962 ( n30492 , n20025 , n8035 );
    not g5963 ( n2656 , n9336 );
    not g5964 ( n9333 , n4160 );
    and g5965 ( n22076 , n31382 , n15328 );
    xnor g5966 ( n23784 , n12071 , n7797 );
    buf g5967 ( n6372 , n9566 );
    not g5968 ( n1367 , n15310 );
    or g5969 ( n21347 , n16048 , n9023 );
    not g5970 ( n27613 , n19916 );
    and g5971 ( n30870 , n27596 , n15614 );
    xnor g5972 ( n3642 , n8766 , n28847 );
    or g5973 ( n12982 , n21612 , n30013 );
    or g5974 ( n16883 , n15736 , n7053 );
    xnor g5975 ( n1876 , n3144 , n8616 );
    xnor g5976 ( n11873 , n25794 , n3810 );
    or g5977 ( n26215 , n12229 , n4241 );
    xor g5978 ( n28611 , n8179 , n6131 );
    and g5979 ( n19031 , n30573 , n13379 );
    or g5980 ( n28030 , n15732 , n16539 );
    xnor g5981 ( n31337 , n6990 , n21577 );
    or g5982 ( n5547 , n5213 , n31522 );
    not g5983 ( n29274 , n3864 );
    not g5984 ( n23762 , n9734 );
    or g5985 ( n26722 , n21604 , n27116 );
    xnor g5986 ( n29844 , n12085 , n14118 );
    xnor g5987 ( n7637 , n29613 , n24067 );
    not g5988 ( n8647 , n8980 );
    xnor g5989 ( n730 , n13974 , n2908 );
    or g5990 ( n18950 , n20987 , n18100 );
    or g5991 ( n15844 , n30096 , n26202 );
    or g5992 ( n4564 , n30212 , n12457 );
    or g5993 ( n30382 , n16194 , n9260 );
    and g5994 ( n3001 , n2606 , n6331 );
    not g5995 ( n21134 , n8561 );
    xnor g5996 ( n14609 , n18671 , n5659 );
    xnor g5997 ( n25807 , n5895 , n6626 );
    xnor g5998 ( n8639 , n2283 , n6018 );
    xnor g5999 ( n3769 , n30673 , n4641 );
    or g6000 ( n28967 , n2136 , n13641 );
    and g6001 ( n5179 , n4269 , n6930 );
    xnor g6002 ( n9341 , n31729 , n11581 );
    not g6003 ( n29855 , n9375 );
    xnor g6004 ( n17385 , n30754 , n28951 );
    and g6005 ( n11734 , n23967 , n2370 );
    not g6006 ( n22299 , n5904 );
    xnor g6007 ( n11714 , n28076 , n1967 );
    nor g6008 ( n28496 , n16135 , n13475 );
    or g6009 ( n31137 , n19078 , n26428 );
    xnor g6010 ( n24526 , n15564 , n23174 );
    xnor g6011 ( n9499 , n15755 , n7799 );
    nor g6012 ( n18754 , n20168 , n1703 );
    not g6013 ( n23344 , n20828 );
    nor g6014 ( n1740 , n18517 , n13232 );
    nor g6015 ( n12148 , n19405 , n28202 );
    xnor g6016 ( n2530 , n6069 , n25182 );
    or g6017 ( n17785 , n4550 , n10512 );
    xnor g6018 ( n26684 , n20802 , n6261 );
    or g6019 ( n7725 , n24136 , n21154 );
    not g6020 ( n26989 , n3642 );
    nor g6021 ( n5337 , n18827 , n29476 );
    nor g6022 ( n26643 , n20038 , n12912 );
    not g6023 ( n13686 , n15612 );
    and g6024 ( n13774 , n30682 , n782 );
    and g6025 ( n31775 , n8502 , n26875 );
    not g6026 ( n25688 , n12335 );
    not g6027 ( n20319 , n30678 );
    not g6028 ( n4316 , n1487 );
    xnor g6029 ( n25724 , n17608 , n14085 );
    and g6030 ( n10025 , n10833 , n19739 );
    xnor g6031 ( n12948 , n17005 , n17090 );
    and g6032 ( n27446 , n10233 , n25582 );
    and g6033 ( n5421 , n26003 , n13126 );
    xor g6034 ( n19570 , n723 , n3571 );
    xnor g6035 ( n1489 , n25126 , n2373 );
    xnor g6036 ( n24463 , n7309 , n5515 );
    not g6037 ( n30552 , n10521 );
    xnor g6038 ( n20735 , n27536 , n28724 );
    not g6039 ( n23633 , n21151 );
    not g6040 ( n6300 , n25462 );
    xnor g6041 ( n14129 , n24151 , n27966 );
    or g6042 ( n19049 , n21853 , n2733 );
    and g6043 ( n4888 , n1758 , n5844 );
    or g6044 ( n4049 , n18452 , n3465 );
    or g6045 ( n29935 , n26968 , n3723 );
    xor g6046 ( n13519 , n23826 , n23959 );
    or g6047 ( n23113 , n23674 , n194 );
    not g6048 ( n24653 , n20486 );
    xnor g6049 ( n11367 , n6527 , n11601 );
    and g6050 ( n14790 , n11821 , n15171 );
    or g6051 ( n10326 , n13700 , n2656 );
    or g6052 ( n15701 , n23362 , n12358 );
    and g6053 ( n8451 , n27242 , n14136 );
    not g6054 ( n6402 , n9759 );
    xnor g6055 ( n10927 , n31895 , n15291 );
    xor g6056 ( n1965 , n7239 , n584 );
    and g6057 ( n27828 , n3020 , n14059 );
    or g6058 ( n27626 , n26204 , n4883 );
    not g6059 ( n16909 , n10289 );
    nor g6060 ( n31432 , n22736 , n5474 );
    or g6061 ( n17991 , n26192 , n10223 );
    or g6062 ( n13339 , n10114 , n23893 );
    nor g6063 ( n17658 , n11665 , n18282 );
    nor g6064 ( n25890 , n6820 , n2596 );
    not g6065 ( n6643 , n7558 );
    not g6066 ( n1516 , n24725 );
    xnor g6067 ( n19587 , n19017 , n23419 );
    or g6068 ( n28382 , n14153 , n24318 );
    xnor g6069 ( n29450 , n25231 , n2631 );
    xnor g6070 ( n1954 , n4166 , n17575 );
    xnor g6071 ( n13505 , n20126 , n9323 );
    or g6072 ( n200 , n31518 , n17925 );
    not g6073 ( n29796 , n25300 );
    not g6074 ( n23873 , n10355 );
    or g6075 ( n18083 , n19567 , n23785 );
    xnor g6076 ( n31445 , n5301 , n18670 );
    nor g6077 ( n11813 , n14235 , n6927 );
    or g6078 ( n15815 , n31487 , n10351 );
    and g6079 ( n27386 , n8873 , n4393 );
    or g6080 ( n13517 , n10552 , n26912 );
    not g6081 ( n10742 , n2681 );
    and g6082 ( n19491 , n16235 , n999 );
    xnor g6083 ( n13450 , n32030 , n5686 );
    or g6084 ( n20673 , n21152 , n17077 );
    xnor g6085 ( n26971 , n28349 , n13565 );
    nor g6086 ( n31949 , n30838 , n7163 );
    xnor g6087 ( n4925 , n12910 , n31470 );
    or g6088 ( n27038 , n15968 , n3660 );
    xnor g6089 ( n2709 , n10710 , n25326 );
    not g6090 ( n12757 , n26102 );
    or g6091 ( n30738 , n4632 , n27205 );
    and g6092 ( n29374 , n25834 , n5324 );
    not g6093 ( n3613 , n22392 );
    and g6094 ( n2793 , n10096 , n3324 );
    xnor g6095 ( n27081 , n8972 , n31728 );
    or g6096 ( n25021 , n21589 , n31864 );
    not g6097 ( n16234 , n7995 );
    or g6098 ( n22008 , n12803 , n1057 );
    and g6099 ( n17551 , n9994 , n5109 );
    not g6100 ( n4914 , n5452 );
    xnor g6101 ( n29078 , n6425 , n27884 );
    xnor g6102 ( n31305 , n3639 , n25699 );
    not g6103 ( n7939 , n28800 );
    and g6104 ( n8616 , n22821 , n22741 );
    or g6105 ( n2598 , n22331 , n7234 );
    and g6106 ( n7263 , n7602 , n15063 );
    or g6107 ( n3929 , n28734 , n31116 );
    buf g6108 ( n10574 , n29919 );
    xnor g6109 ( n23591 , n31766 , n5701 );
    not g6110 ( n20141 , n13186 );
    and g6111 ( n8467 , n266 , n31827 );
    or g6112 ( n27017 , n1153 , n7977 );
    not g6113 ( n11970 , n21156 );
    and g6114 ( n9001 , n17516 , n15053 );
    not g6115 ( n25305 , n445 );
    or g6116 ( n13036 , n17779 , n30599 );
    xnor g6117 ( n27469 , n11063 , n18753 );
    and g6118 ( n28313 , n12883 , n10053 );
    and g6119 ( n3275 , n1624 , n16818 );
    not g6120 ( n15716 , n18040 );
    not g6121 ( n7720 , n21487 );
    and g6122 ( n17187 , n5785 , n16904 );
    not g6123 ( n13782 , n30541 );
    not g6124 ( n16690 , n17647 );
    or g6125 ( n28959 , n31965 , n10980 );
    not g6126 ( n1006 , n19231 );
    xnor g6127 ( n25386 , n17197 , n10040 );
    and g6128 ( n17164 , n16684 , n9915 );
    xnor g6129 ( n15904 , n1207 , n19680 );
    xnor g6130 ( n1545 , n30857 , n303 );
    or g6131 ( n28812 , n6842 , n13771 );
    or g6132 ( n31223 , n7180 , n16134 );
    nor g6133 ( n11925 , n20038 , n25587 );
    and g6134 ( n866 , n12923 , n5678 );
    and g6135 ( n4798 , n10892 , n13847 );
    or g6136 ( n3238 , n31469 , n446 );
    nor g6137 ( n29030 , n24484 , n24672 );
    not g6138 ( n27091 , n22708 );
    not g6139 ( n10729 , n10460 );
    or g6140 ( n14389 , n30356 , n319 );
    or g6141 ( n5486 , n9886 , n1940 );
    not g6142 ( n8311 , n3773 );
    and g6143 ( n7803 , n9923 , n16352 );
    or g6144 ( n29555 , n25890 , n25560 );
    or g6145 ( n16999 , n12928 , n24625 );
    xnor g6146 ( n24581 , n22886 , n2610 );
    not g6147 ( n11916 , n5388 );
    not g6148 ( n23726 , n21960 );
    or g6149 ( n5219 , n4599 , n29332 );
    xnor g6150 ( n24795 , n10143 , n19099 );
    xnor g6151 ( n22828 , n25384 , n6338 );
    nor g6152 ( n4576 , n10643 , n14875 );
    or g6153 ( n10284 , n24627 , n26872 );
    not g6154 ( n23082 , n14013 );
    or g6155 ( n16245 , n3407 , n18367 );
    or g6156 ( n19446 , n28033 , n7331 );
    xnor g6157 ( n23798 , n26786 , n6141 );
    or g6158 ( n22190 , n4409 , n4894 );
    xnor g6159 ( n6727 , n28217 , n848 );
    not g6160 ( n18227 , n20747 );
    and g6161 ( n639 , n3957 , n4291 );
    not g6162 ( n23618 , n25336 );
    nor g6163 ( n29460 , n23669 , n6371 );
    not g6164 ( n26748 , n22422 );
    nor g6165 ( n30034 , n15301 , n11355 );
    or g6166 ( n15859 , n5690 , n19410 );
    xnor g6167 ( n7969 , n31785 , n19508 );
    not g6168 ( n8507 , n27199 );
    or g6169 ( n20928 , n15717 , n20596 );
    not g6170 ( n1952 , n5427 );
    xnor g6171 ( n17955 , n3782 , n3907 );
    xnor g6172 ( n1908 , n23146 , n5099 );
    xnor g6173 ( n6942 , n20572 , n8705 );
    xnor g6174 ( n31221 , n22670 , n14979 );
    not g6175 ( n9187 , n21648 );
    or g6176 ( n1452 , n20396 , n30621 );
    and g6177 ( n26897 , n5491 , n30711 );
    not g6178 ( n8211 , n26620 );
    nor g6179 ( n24485 , n18229 , n22842 );
    not g6180 ( n27013 , n26176 );
    nor g6181 ( n25430 , n25527 , n12602 );
    not g6182 ( n1521 , n13286 );
    or g6183 ( n21149 , n25686 , n2344 );
    or g6184 ( n2305 , n2555 , n25563 );
    or g6185 ( n29617 , n26831 , n25483 );
    not g6186 ( n20789 , n6579 );
    not g6187 ( n19344 , n12685 );
    xnor g6188 ( n983 , n11640 , n15999 );
    and g6189 ( n29821 , n25669 , n21493 );
    or g6190 ( n17850 , n1285 , n14376 );
    nor g6191 ( n17327 , n16075 , n14106 );
    xnor g6192 ( n13642 , n27126 , n3312 );
    and g6193 ( n112 , n8010 , n25449 );
    nor g6194 ( n24090 , n20313 , n11305 );
    not g6195 ( n21525 , n4901 );
    not g6196 ( n30635 , n24518 );
    not g6197 ( n6446 , n11701 );
    or g6198 ( n26272 , n14030 , n14755 );
    not g6199 ( n24889 , n21909 );
    xnor g6200 ( n4742 , n13303 , n3006 );
    and g6201 ( n19611 , n25724 , n5503 );
    or g6202 ( n23959 , n11692 , n8435 );
    not g6203 ( n23931 , n13836 );
    and g6204 ( n21838 , n20426 , n20048 );
    not g6205 ( n2653 , n29604 );
    and g6206 ( n16989 , n2342 , n9651 );
    buf g6207 ( n667 , n28763 );
    not g6208 ( n20208 , n6578 );
    and g6209 ( n16777 , n10789 , n8703 );
    or g6210 ( n11890 , n22709 , n12534 );
    xor g6211 ( n6735 , n18560 , n26435 );
    not g6212 ( n22044 , n16617 );
    xor g6213 ( n24003 , n7652 , n13689 );
    xnor g6214 ( n18629 , n20223 , n26518 );
    and g6215 ( n15089 , n25038 , n11170 );
    or g6216 ( n5617 , n23539 , n12150 );
    xnor g6217 ( n29364 , n26675 , n29447 );
    not g6218 ( n31446 , n5839 );
    not g6219 ( n27589 , n13682 );
    or g6220 ( n17055 , n9646 , n24611 );
    and g6221 ( n22639 , n27225 , n9083 );
    and g6222 ( n21798 , n9962 , n19217 );
    or g6223 ( n29268 , n30836 , n23717 );
    xnor g6224 ( n19337 , n22053 , n14558 );
    not g6225 ( n1600 , n11736 );
    nor g6226 ( n29068 , n17356 , n15083 );
    not g6227 ( n4474 , n22690 );
    xnor g6228 ( n12160 , n29609 , n10163 );
    and g6229 ( n30251 , n31709 , n5089 );
    or g6230 ( n24041 , n28921 , n10313 );
    not g6231 ( n6047 , n31461 );
    and g6232 ( n27953 , n7653 , n7211 );
    nor g6233 ( n14033 , n16815 , n3377 );
    and g6234 ( n11149 , n29603 , n17395 );
    xnor g6235 ( n24083 , n9639 , n21137 );
    not g6236 ( n18807 , n8228 );
    nor g6237 ( n5068 , n3051 , n25116 );
    xnor g6238 ( n23558 , n28138 , n29412 );
    and g6239 ( n7982 , n8165 , n12491 );
    or g6240 ( n25820 , n3123 , n2515 );
    xnor g6241 ( n20563 , n508 , n8321 );
    not g6242 ( n13889 , n24355 );
    not g6243 ( n30597 , n19805 );
    not g6244 ( n16322 , n3993 );
    xnor g6245 ( n13565 , n28560 , n14858 );
    and g6246 ( n10901 , n9188 , n25323 );
    xnor g6247 ( n24321 , n23365 , n18380 );
    xnor g6248 ( n30625 , n5524 , n8715 );
    or g6249 ( n14217 , n7473 , n17071 );
    xnor g6250 ( n5637 , n19905 , n16578 );
    xnor g6251 ( n10255 , n17096 , n25825 );
    or g6252 ( n25683 , n19524 , n4960 );
    or g6253 ( n23580 , n10942 , n1355 );
    or g6254 ( n9027 , n17090 , n22088 );
    and g6255 ( n19788 , n20429 , n22430 );
    and g6256 ( n3714 , n20537 , n20884 );
    xnor g6257 ( n28404 , n16943 , n6388 );
    or g6258 ( n9741 , n12490 , n12755 );
    not g6259 ( n29676 , n6755 );
    or g6260 ( n22599 , n6355 , n1844 );
    and g6261 ( n8693 , n22407 , n30983 );
    and g6262 ( n31472 , n1323 , n12303 );
    xnor g6263 ( n15618 , n6618 , n24974 );
    xnor g6264 ( n734 , n2051 , n5203 );
    and g6265 ( n28266 , n18801 , n30243 );
    and g6266 ( n11474 , n30938 , n4049 );
    xnor g6267 ( n14583 , n7086 , n23232 );
    xnor g6268 ( n11161 , n23960 , n2934 );
    not g6269 ( n21582 , n25746 );
    and g6270 ( n25739 , n5260 , n11060 );
    or g6271 ( n7616 , n23247 , n1683 );
    xnor g6272 ( n18890 , n26974 , n10676 );
    or g6273 ( n6028 , n12542 , n2014 );
    and g6274 ( n20700 , n28881 , n9356 );
    not g6275 ( n7980 , n4628 );
    and g6276 ( n28246 , n11772 , n12134 );
    xnor g6277 ( n27900 , n22198 , n1745 );
    or g6278 ( n9403 , n23195 , n7957 );
    and g6279 ( n3564 , n1605 , n5303 );
    not g6280 ( n21141 , n21063 );
    or g6281 ( n31279 , n1380 , n5992 );
    not g6282 ( n27605 , n19566 );
    not g6283 ( n7258 , n31165 );
    not g6284 ( n29552 , n12803 );
    or g6285 ( n1009 , n22922 , n19300 );
    or g6286 ( n25263 , n5375 , n31956 );
    not g6287 ( n17218 , n6012 );
    xnor g6288 ( n18417 , n22800 , n20319 );
    nor g6289 ( n30485 , n11610 , n7669 );
    xnor g6290 ( n17108 , n10078 , n26878 );
    xnor g6291 ( n26603 , n20588 , n14864 );
    or g6292 ( n12643 , n14525 , n28414 );
    xnor g6293 ( n16826 , n2761 , n13551 );
    xnor g6294 ( n296 , n16481 , n16651 );
    nor g6295 ( n7744 , n12796 , n16809 );
    xnor g6296 ( n28497 , n24782 , n25001 );
    or g6297 ( n13627 , n11867 , n26745 );
    xnor g6298 ( n1043 , n1742 , n31727 );
    or g6299 ( n27171 , n9763 , n16083 );
    nor g6300 ( n28301 , n19651 , n22123 );
    not g6301 ( n26632 , n24235 );
    or g6302 ( n3049 , n8901 , n20013 );
    or g6303 ( n10874 , n11684 , n11501 );
    and g6304 ( n22890 , n12655 , n9431 );
    not g6305 ( n17093 , n24070 );
    nor g6306 ( n16495 , n213 , n11284 );
    not g6307 ( n18229 , n9691 );
    not g6308 ( n30194 , n16476 );
    or g6309 ( n3860 , n347 , n24190 );
    xnor g6310 ( n20434 , n23675 , n11109 );
    or g6311 ( n20307 , n27893 , n4520 );
    or g6312 ( n3969 , n14625 , n17658 );
    or g6313 ( n31114 , n14675 , n16466 );
    or g6314 ( n6202 , n24040 , n13587 );
    not g6315 ( n30057 , n26859 );
    or g6316 ( n27846 , n4394 , n6035 );
    xnor g6317 ( n10296 , n9231 , n20494 );
    xnor g6318 ( n21973 , n12829 , n23976 );
    or g6319 ( n21913 , n18802 , n26146 );
    xnor g6320 ( n31539 , n28273 , n6574 );
    or g6321 ( n22668 , n6861 , n21663 );
    xnor g6322 ( n19904 , n26082 , n6957 );
    not g6323 ( n11097 , n15531 );
    xnor g6324 ( n21694 , n850 , n15414 );
    and g6325 ( n5394 , n28385 , n17813 );
    not g6326 ( n30232 , n22154 );
    not g6327 ( n8392 , n3531 );
    xnor g6328 ( n17053 , n12181 , n25242 );
    nor g6329 ( n28355 , n23772 , n3743 );
    and g6330 ( n12532 , n24117 , n22444 );
    not g6331 ( n21820 , n24422 );
    not g6332 ( n11103 , n31761 );
    and g6333 ( n3344 , n24565 , n10161 );
    not g6334 ( n8266 , n28695 );
    not g6335 ( n9312 , n3591 );
    or g6336 ( n13593 , n9744 , n15010 );
    not g6337 ( n18746 , n30514 );
    not g6338 ( n27936 , n17255 );
    and g6339 ( n2992 , n9332 , n27323 );
    nor g6340 ( n6964 , n27227 , n11110 );
    not g6341 ( n4872 , n6465 );
    not g6342 ( n10431 , n6391 );
    nor g6343 ( n4282 , n6172 , n20510 );
    nor g6344 ( n4019 , n30534 , n12282 );
    not g6345 ( n10658 , n3108 );
    or g6346 ( n9379 , n15733 , n7812 );
    and g6347 ( n10843 , n2893 , n14948 );
    xnor g6348 ( n12798 , n27455 , n2477 );
    nor g6349 ( n2237 , n18210 , n17898 );
    nor g6350 ( n19742 , n27443 , n4848 );
    not g6351 ( n713 , n9280 );
    or g6352 ( n24686 , n28149 , n31031 );
    or g6353 ( n15740 , n1123 , n16988 );
    and g6354 ( n28577 , n29409 , n29184 );
    not g6355 ( n3010 , n19476 );
    not g6356 ( n14574 , n220 );
    not g6357 ( n4707 , n19651 );
    xnor g6358 ( n11937 , n10985 , n10574 );
    nor g6359 ( n19936 , n19538 , n3057 );
    or g6360 ( n2257 , n14783 , n28516 );
    or g6361 ( n23822 , n17021 , n29564 );
    or g6362 ( n19072 , n27765 , n7259 );
    not g6363 ( n5248 , n17379 );
    or g6364 ( n25160 , n10668 , n20879 );
    or g6365 ( n665 , n26043 , n26567 );
    and g6366 ( n13942 , n31418 , n7322 );
    and g6367 ( n17198 , n5681 , n16976 );
    or g6368 ( n7521 , n20187 , n9269 );
    or g6369 ( n27869 , n17 , n13986 );
    and g6370 ( n28101 , n24718 , n17152 );
    or g6371 ( n24403 , n9855 , n12581 );
    and g6372 ( n5750 , n15364 , n18241 );
    and g6373 ( n23413 , n25160 , n3328 );
    nor g6374 ( n15140 , n9097 , n8945 );
    xnor g6375 ( n30231 , n4944 , n10546 );
    xnor g6376 ( n7780 , n31537 , n15542 );
    or g6377 ( n18579 , n10062 , n1682 );
    xnor g6378 ( n12896 , n14074 , n16299 );
    not g6379 ( n21173 , n8919 );
    xnor g6380 ( n3494 , n7857 , n19300 );
    not g6381 ( n5276 , n21921 );
    or g6382 ( n3609 , n12485 , n28544 );
    and g6383 ( n22967 , n26921 , n601 );
    not g6384 ( n30820 , n7409 );
    and g6385 ( n5913 , n6190 , n23631 );
    or g6386 ( n15212 , n2548 , n31090 );
    or g6387 ( n27835 , n7727 , n1106 );
    and g6388 ( n31092 , n16575 , n11641 );
    not g6389 ( n24969 , n28180 );
    or g6390 ( n13511 , n17669 , n5899 );
    and g6391 ( n18054 , n21663 , n24614 );
    xnor g6392 ( n10705 , n16800 , n19405 );
    not g6393 ( n20720 , n15417 );
    not g6394 ( n6720 , n30062 );
    xnor g6395 ( n10118 , n18250 , n18648 );
    nor g6396 ( n26840 , n3405 , n7982 );
    xnor g6397 ( n13345 , n31347 , n25432 );
    not g6398 ( n3948 , n15791 );
    or g6399 ( n12957 , n23145 , n13516 );
    not g6400 ( n21654 , n752 );
    and g6401 ( n2977 , n25780 , n31724 );
    or g6402 ( n20668 , n3 , n25354 );
    and g6403 ( n19531 , n25030 , n29139 );
    xnor g6404 ( n19474 , n20733 , n4495 );
    xnor g6405 ( n13397 , n1187 , n17122 );
    not g6406 ( n7283 , n3661 );
    or g6407 ( n27870 , n18443 , n6992 );
    and g6408 ( n18122 , n9552 , n15005 );
    not g6409 ( n24095 , n7658 );
    or g6410 ( n29916 , n15272 , n9531 );
    not g6411 ( n26131 , n14288 );
    not g6412 ( n18681 , n7549 );
    not g6413 ( n25091 , n7444 );
    or g6414 ( n28501 , n4393 , n23160 );
    xnor g6415 ( n15501 , n6377 , n2200 );
    or g6416 ( n22175 , n4974 , n27173 );
    xor g6417 ( n25247 , n11109 , n3816 );
    or g6418 ( n556 , n27776 , n9186 );
    xnor g6419 ( n24946 , n3236 , n11940 );
    xnor g6420 ( n18140 , n14844 , n717 );
    not g6421 ( n6633 , n223 );
    or g6422 ( n14146 , n26286 , n29207 );
    xnor g6423 ( n18654 , n19827 , n15040 );
    not g6424 ( n24287 , n30904 );
    and g6425 ( n23527 , n8403 , n15588 );
    nor g6426 ( n21086 , n3863 , n10047 );
    not g6427 ( n16576 , n21295 );
    not g6428 ( n20310 , n18596 );
    nor g6429 ( n5346 , n31106 , n24792 );
    xnor g6430 ( n12821 , n14784 , n29795 );
    or g6431 ( n8210 , n8539 , n10530 );
    or g6432 ( n13069 , n22963 , n28480 );
    and g6433 ( n4181 , n21403 , n24248 );
    xor g6434 ( n14209 , n1312 , n13712 );
    not g6435 ( n27316 , n24694 );
    xnor g6436 ( n17199 , n26191 , n22512 );
    nor g6437 ( n21162 , n28375 , n9711 );
    xnor g6438 ( n17880 , n16037 , n10048 );
    xnor g6439 ( n800 , n22461 , n6469 );
    or g6440 ( n31063 , n2740 , n13782 );
    xnor g6441 ( n13298 , n1797 , n30005 );
    and g6442 ( n29954 , n24397 , n9428 );
    not g6443 ( n26464 , n26707 );
    not g6444 ( n18063 , n17798 );
    and g6445 ( n5956 , n12170 , n17227 );
    not g6446 ( n9793 , n1718 );
    not g6447 ( n17299 , n25395 );
    xnor g6448 ( n817 , n20796 , n5560 );
    nor g6449 ( n29047 , n3034 , n23810 );
    or g6450 ( n3852 , n31123 , n30750 );
    or g6451 ( n12177 , n21660 , n2586 );
    not g6452 ( n23850 , n10639 );
    not g6453 ( n8052 , n4751 );
    xnor g6454 ( n21408 , n27738 , n3513 );
    or g6455 ( n15157 , n22675 , n1424 );
    xnor g6456 ( n5703 , n13725 , n8834 );
    or g6457 ( n5534 , n6329 , n20219 );
    and g6458 ( n30673 , n26042 , n17827 );
    xnor g6459 ( n7272 , n28013 , n31711 );
    or g6460 ( n8408 , n9695 , n24925 );
    not g6461 ( n1278 , n19331 );
    xnor g6462 ( n1539 , n2785 , n18884 );
    nor g6463 ( n3838 , n15573 , n9798 );
    nor g6464 ( n22143 , n16778 , n29288 );
    not g6465 ( n27860 , n727 );
    or g6466 ( n29767 , n20829 , n9393 );
    xnor g6467 ( n12689 , n952 , n21114 );
    or g6468 ( n15773 , n29373 , n11144 );
    not g6469 ( n17076 , n16409 );
    xnor g6470 ( n1951 , n3688 , n2934 );
    xnor g6471 ( n23578 , n9488 , n8804 );
    xnor g6472 ( n25211 , n3863 , n21508 );
    not g6473 ( n22660 , n5726 );
    xnor g6474 ( n14641 , n27300 , n18755 );
    not g6475 ( n20705 , n15109 );
    xnor g6476 ( n25661 , n17771 , n7655 );
    xor g6477 ( n15112 , n17533 , n4662 );
    or g6478 ( n18569 , n13916 , n2850 );
    and g6479 ( n28498 , n11509 , n11650 );
    nor g6480 ( n20539 , n3259 , n2883 );
    or g6481 ( n5698 , n30398 , n11874 );
    xnor g6482 ( n6642 , n19073 , n15340 );
    not g6483 ( n392 , n1342 );
    xnor g6484 ( n7852 , n17148 , n28345 );
    not g6485 ( n6955 , n30828 );
    or g6486 ( n17984 , n7445 , n8734 );
    xnor g6487 ( n5907 , n30442 , n20006 );
    or g6488 ( n30147 , n12661 , n21550 );
    nor g6489 ( n13678 , n2021 , n25198 );
    or g6490 ( n885 , n15173 , n25153 );
    and g6491 ( n31841 , n15383 , n16745 );
    or g6492 ( n9420 , n30025 , n23090 );
    and g6493 ( n10381 , n25055 , n26811 );
    not g6494 ( n31160 , n11045 );
    or g6495 ( n29099 , n31342 , n6892 );
    nor g6496 ( n26257 , n31595 , n15797 );
    not g6497 ( n23932 , n2798 );
    and g6498 ( n30328 , n5983 , n21428 );
    xnor g6499 ( n22388 , n2819 , n29337 );
    xnor g6500 ( n12297 , n23620 , n14828 );
    xnor g6501 ( n29984 , n13757 , n3346 );
    and g6502 ( n29685 , n26374 , n12607 );
    and g6503 ( n22859 , n3609 , n24346 );
    and g6504 ( n17241 , n17826 , n29471 );
    not g6505 ( n12624 , n26321 );
    and g6506 ( n18457 , n10763 , n27710 );
    and g6507 ( n28434 , n4902 , n1003 );
    and g6508 ( n31934 , n7789 , n5923 );
    and g6509 ( n29773 , n28224 , n15990 );
    xnor g6510 ( n9155 , n3145 , n8200 );
    xnor g6511 ( n12216 , n12097 , n23804 );
    xnor g6512 ( n24144 , n16097 , n30800 );
    not g6513 ( n5287 , n29903 );
    xnor g6514 ( n8076 , n15485 , n23248 );
    not g6515 ( n25007 , n18237 );
    xnor g6516 ( n26963 , n19448 , n12136 );
    xnor g6517 ( n27636 , n8743 , n18904 );
    not g6518 ( n7025 , n30476 );
    not g6519 ( n1573 , n30412 );
    not g6520 ( n29987 , n16350 );
    and g6521 ( n31874 , n3201 , n4693 );
    and g6522 ( n4940 , n28861 , n23055 );
    xnor g6523 ( n12877 , n17321 , n23145 );
    and g6524 ( n29531 , n15114 , n8362 );
    not g6525 ( n5906 , n31481 );
    or g6526 ( n10481 , n21681 , n23827 );
    not g6527 ( n14534 , n459 );
    or g6528 ( n8752 , n26841 , n438 );
    xnor g6529 ( n22667 , n14453 , n20724 );
    xnor g6530 ( n10250 , n16200 , n3688 );
    xor g6531 ( n15609 , n27766 , n21515 );
    and g6532 ( n24088 , n19569 , n31896 );
    or g6533 ( n14251 , n30521 , n9932 );
    xnor g6534 ( n1180 , n19138 , n15266 );
    not g6535 ( n17480 , n28678 );
    xnor g6536 ( n600 , n1688 , n24148 );
    or g6537 ( n31529 , n1093 , n2241 );
    not g6538 ( n5622 , n21159 );
    xnor g6539 ( n14598 , n30376 , n26056 );
    and g6540 ( n14329 , n5873 , n5150 );
    not g6541 ( n17100 , n19120 );
    or g6542 ( n26645 , n28770 , n8308 );
    not g6543 ( n21342 , n31928 );
    xnor g6544 ( n3249 , n6686 , n1177 );
    not g6545 ( n4410 , n5328 );
    nor g6546 ( n26420 , n12859 , n5973 );
    xnor g6547 ( n5813 , n25866 , n23635 );
    or g6548 ( n27749 , n12396 , n28403 );
    xnor g6549 ( n20866 , n22082 , n7656 );
    xnor g6550 ( n14630 , n14017 , n20845 );
    not g6551 ( n12157 , n11742 );
    or g6552 ( n27194 , n8528 , n14845 );
    not g6553 ( n21831 , n8760 );
    or g6554 ( n314 , n20254 , n31511 );
    xnor g6555 ( n16321 , n15384 , n23491 );
    xnor g6556 ( n23514 , n13536 , n9638 );
    nor g6557 ( n24932 , n15724 , n20575 );
    or g6558 ( n17020 , n19955 , n15867 );
    nor g6559 ( n14721 , n16831 , n19250 );
    nor g6560 ( n22709 , n27131 , n1877 );
    or g6561 ( n26575 , n31229 , n22565 );
    and g6562 ( n30766 , n21035 , n19503 );
    or g6563 ( n8962 , n11746 , n20425 );
    xnor g6564 ( n20418 , n3680 , n25889 );
    buf g6565 ( n19590 , n25718 );
    nor g6566 ( n5660 , n29153 , n4612 );
    not g6567 ( n10515 , n9391 );
    and g6568 ( n25573 , n29405 , n8904 );
    not g6569 ( n20834 , n26300 );
    or g6570 ( n27800 , n30666 , n28834 );
    not g6571 ( n4906 , n28724 );
    nor g6572 ( n14884 , n31813 , n14069 );
    and g6573 ( n8349 , n19402 , n16118 );
    not g6574 ( n2416 , n11192 );
    and g6575 ( n3805 , n15483 , n9166 );
    or g6576 ( n1138 , n27583 , n17365 );
    or g6577 ( n585 , n2939 , n12514 );
    xnor g6578 ( n29421 , n5983 , n9037 );
    xnor g6579 ( n31433 , n1535 , n19221 );
    not g6580 ( n7598 , n27602 );
    not g6581 ( n8003 , n212 );
    or g6582 ( n7561 , n29975 , n26853 );
    and g6583 ( n17680 , n12302 , n10987 );
    not g6584 ( n17928 , n31320 );
    not g6585 ( n18709 , n20692 );
    and g6586 ( n23946 , n9441 , n15214 );
    and g6587 ( n1523 , n23737 , n30725 );
    not g6588 ( n14798 , n16478 );
    or g6589 ( n9218 , n6653 , n9486 );
    and g6590 ( n15781 , n2880 , n19365 );
    not g6591 ( n22493 , n7414 );
    and g6592 ( n30237 , n20162 , n20102 );
    or g6593 ( n18081 , n19223 , n28353 );
    not g6594 ( n13704 , n9650 );
    nor g6595 ( n6405 , n22423 , n12035 );
    xnor g6596 ( n10514 , n23827 , n24224 );
    xnor g6597 ( n8702 , n24594 , n12117 );
    not g6598 ( n26888 , n3189 );
    and g6599 ( n22206 , n9057 , n9572 );
    not g6600 ( n17670 , n15085 );
    not g6601 ( n28934 , n30957 );
    or g6602 ( n11871 , n4525 , n19803 );
    xnor g6603 ( n29832 , n227 , n19572 );
    xnor g6604 ( n10232 , n29794 , n4924 );
    and g6605 ( n1340 , n18354 , n21053 );
    or g6606 ( n10341 , n1359 , n19605 );
    or g6607 ( n5632 , n13113 , n21468 );
    xnor g6608 ( n13858 , n5301 , n29830 );
    xnor g6609 ( n22921 , n23873 , n5105 );
    or g6610 ( n22822 , n3663 , n14170 );
    and g6611 ( n12167 , n23591 , n10043 );
    and g6612 ( n19409 , n16569 , n21607 );
    xnor g6613 ( n12858 , n24351 , n13528 );
    xnor g6614 ( n29725 , n16531 , n1195 );
    not g6615 ( n14133 , n11601 );
    nor g6616 ( n19362 , n31168 , n16890 );
    not g6617 ( n20643 , n11975 );
    and g6618 ( n7667 , n18692 , n6252 );
    xnor g6619 ( n21303 , n18798 , n22449 );
    or g6620 ( n24870 , n1963 , n7667 );
    not g6621 ( n31912 , n1368 );
    not g6622 ( n20765 , n6527 );
    or g6623 ( n2896 , n25849 , n14726 );
    xnor g6624 ( n30455 , n21390 , n29444 );
    xnor g6625 ( n1837 , n9773 , n26467 );
    or g6626 ( n1556 , n729 , n21713 );
    and g6627 ( n6081 , n3114 , n18144 );
    or g6628 ( n8027 , n24006 , n8471 );
    not g6629 ( n19641 , n17227 );
    not g6630 ( n29751 , n3240 );
    not g6631 ( n25373 , n28237 );
    and g6632 ( n19112 , n31569 , n26134 );
    or g6633 ( n18205 , n21093 , n15703 );
    or g6634 ( n16172 , n30139 , n14700 );
    or g6635 ( n2445 , n6275 , n12406 );
    not g6636 ( n21919 , n24773 );
    and g6637 ( n13916 , n7957 , n23195 );
    and g6638 ( n8342 , n24947 , n5473 );
    not g6639 ( n4767 , n4175 );
    not g6640 ( n31646 , n4956 );
    nor g6641 ( n18938 , n26558 , n5221 );
    or g6642 ( n24430 , n24579 , n3158 );
    not g6643 ( n12315 , n2938 );
    or g6644 ( n25323 , n21849 , n25971 );
    or g6645 ( n24635 , n25003 , n11067 );
    not g6646 ( n9715 , n15300 );
    not g6647 ( n27285 , n18575 );
    or g6648 ( n27802 , n6600 , n13013 );
    nor g6649 ( n26092 , n5265 , n5011 );
    not g6650 ( n29228 , n12777 );
    or g6651 ( n18332 , n393 , n137 );
    not g6652 ( n19808 , n8538 );
    or g6653 ( n1103 , n3145 , n11097 );
    not g6654 ( n6800 , n9325 );
    and g6655 ( n12709 , n14309 , n16614 );
    not g6656 ( n5847 , n30274 );
    not g6657 ( n16756 , n13410 );
    and g6658 ( n20696 , n17303 , n29884 );
    not g6659 ( n29812 , n16333 );
    not g6660 ( n14354 , n15683 );
    or g6661 ( n26382 , n27335 , n12377 );
    or g6662 ( n8441 , n8882 , n5478 );
    nor g6663 ( n24721 , n27731 , n31196 );
    not g6664 ( n8137 , n7109 );
    xnor g6665 ( n6320 , n14621 , n30120 );
    xnor g6666 ( n7212 , n9336 , n13700 );
    xnor g6667 ( n29734 , n3787 , n7655 );
    and g6668 ( n18036 , n20257 , n12132 );
    or g6669 ( n27045 , n15 , n64 );
    xnor g6670 ( n9339 , n28922 , n19799 );
    not g6671 ( n16154 , n541 );
    or g6672 ( n11695 , n27018 , n20112 );
    nor g6673 ( n11703 , n2311 , n25122 );
    not g6674 ( n19577 , n20871 );
    not g6675 ( n19502 , n15357 );
    xnor g6676 ( n24175 , n28097 , n16948 );
    not g6677 ( n15329 , n7988 );
    and g6678 ( n7950 , n7908 , n10431 );
    and g6679 ( n12793 , n25717 , n29532 );
    and g6680 ( n5059 , n13243 , n8834 );
    not g6681 ( n14876 , n2071 );
    and g6682 ( n25560 , n28181 , n7437 );
    and g6683 ( n12934 , n30594 , n3312 );
    and g6684 ( n13792 , n2307 , n18217 );
    or g6685 ( n17937 , n7399 , n30849 );
    and g6686 ( n7481 , n9780 , n22322 );
    nor g6687 ( n3167 , n7705 , n30207 );
    not g6688 ( n20786 , n23270 );
    xor g6689 ( n23044 , n148 , n25285 );
    xnor g6690 ( n10177 , n1802 , n28788 );
    and g6691 ( n23524 , n21860 , n20491 );
    xnor g6692 ( n12360 , n30045 , n10433 );
    or g6693 ( n22785 , n7512 , n13316 );
    and g6694 ( n29442 , n6905 , n9016 );
    not g6695 ( n278 , n26429 );
    or g6696 ( n22017 , n13725 , n1841 );
    not g6697 ( n2464 , n25066 );
    not g6698 ( n1427 , n10558 );
    not g6699 ( n22268 , n1191 );
    and g6700 ( n23123 , n10107 , n30476 );
    nor g6701 ( n1441 , n3244 , n28134 );
    not g6702 ( n25397 , n9152 );
    or g6703 ( n27822 , n8061 , n18269 );
    xnor g6704 ( n27818 , n15462 , n20447 );
    nor g6705 ( n126 , n18548 , n7664 );
    or g6706 ( n10164 , n12616 , n13206 );
    or g6707 ( n22585 , n11636 , n20383 );
    and g6708 ( n15466 , n28310 , n17840 );
    or g6709 ( n26216 , n166 , n13618 );
    not g6710 ( n26544 , n28230 );
    nor g6711 ( n29958 , n24094 , n18695 );
    xnor g6712 ( n2348 , n14531 , n16795 );
    or g6713 ( n5801 , n3091 , n18550 );
    or g6714 ( n1121 , n3812 , n29685 );
    xnor g6715 ( n6630 , n15331 , n31355 );
    xnor g6716 ( n4611 , n8088 , n6281 );
    and g6717 ( n1868 , n27130 , n19135 );
    or g6718 ( n17587 , n3810 , n942 );
    xnor g6719 ( n1792 , n11792 , n27501 );
    nor g6720 ( n27054 , n4571 , n3592 );
    or g6721 ( n19824 , n1941 , n23579 );
    not g6722 ( n26070 , n27271 );
    not g6723 ( n475 , n21229 );
    or g6724 ( n22160 , n17723 , n27425 );
    xnor g6725 ( n18156 , n29103 , n22187 );
    not g6726 ( n26795 , n14458 );
    xnor g6727 ( n2335 , n10490 , n6196 );
    and g6728 ( n18307 , n24154 , n24378 );
    and g6729 ( n20021 , n30976 , n20406 );
    not g6730 ( n25001 , n3678 );
    and g6731 ( n8723 , n29551 , n10906 );
    or g6732 ( n9465 , n9310 , n2315 );
    xnor g6733 ( n29192 , n574 , n5728 );
    or g6734 ( n10654 , n8586 , n21667 );
    not g6735 ( n1828 , n19880 );
    or g6736 ( n26253 , n12253 , n5729 );
    nor g6737 ( n21225 , n6115 , n12258 );
    buf g6738 ( n6370 , n2950 );
    and g6739 ( n14726 , n4616 , n4540 );
    not g6740 ( n13486 , n17724 );
    nor g6741 ( n21411 , n30593 , n20779 );
    and g6742 ( n28974 , n15613 , n21310 );
    not g6743 ( n11344 , n21540 );
    xnor g6744 ( n23108 , n6518 , n21892 );
    not g6745 ( n8273 , n22647 );
    xnor g6746 ( n21187 , n8328 , n11494 );
    or g6747 ( n6225 , n97 , n2150 );
    xnor g6748 ( n1007 , n399 , n25334 );
    not g6749 ( n30069 , n10973 );
    or g6750 ( n21024 , n14874 , n22840 );
    or g6751 ( n29819 , n604 , n16064 );
    not g6752 ( n12403 , n24056 );
    xnor g6753 ( n9303 , n31775 , n2788 );
    and g6754 ( n15929 , n27386 , n24464 );
    or g6755 ( n839 , n15555 , n5663 );
    and g6756 ( n979 , n19324 , n25385 );
    and g6757 ( n13638 , n1475 , n27762 );
    not g6758 ( n2660 , n24066 );
    not g6759 ( n3481 , n26636 );
    and g6760 ( n29570 , n26289 , n6141 );
    and g6761 ( n17598 , n26382 , n12615 );
    and g6762 ( n25101 , n30609 , n16665 );
    not g6763 ( n15624 , n12207 );
    xnor g6764 ( n12347 , n21982 , n24522 );
    not g6765 ( n20014 , n23784 );
    not g6766 ( n10631 , n23270 );
    and g6767 ( n22253 , n41 , n3268 );
    nor g6768 ( n12124 , n9835 , n4004 );
    xnor g6769 ( n1738 , n6960 , n8454 );
    nor g6770 ( n4310 , n3765 , n2963 );
    and g6771 ( n15268 , n6879 , n11608 );
    xnor g6772 ( n17278 , n14333 , n14962 );
    not g6773 ( n5065 , n17010 );
    and g6774 ( n16050 , n20701 , n4685 );
    not g6775 ( n28882 , n24436 );
    and g6776 ( n4262 , n518 , n8834 );
    or g6777 ( n5945 , n21673 , n20639 );
    xnor g6778 ( n22575 , n30215 , n2377 );
    and g6779 ( n25602 , n26574 , n16935 );
    not g6780 ( n21524 , n17930 );
    and g6781 ( n14773 , n29140 , n11584 );
    nor g6782 ( n12616 , n20881 , n14119 );
    or g6783 ( n9513 , n31371 , n28423 );
    and g6784 ( n18494 , n27539 , n17656 );
    and g6785 ( n8257 , n31346 , n25530 );
    xnor g6786 ( n31217 , n23492 , n29387 );
    not g6787 ( n1368 , n16011 );
    xor g6788 ( n292 , n16356 , n8908 );
    not g6789 ( n21714 , n13795 );
    xnor g6790 ( n23060 , n27669 , n20114 );
    xnor g6791 ( n20812 , n23214 , n22120 );
    xnor g6792 ( n6362 , n4613 , n23323 );
    and g6793 ( n25463 , n4921 , n24058 );
    or g6794 ( n28104 , n28926 , n25606 );
    xnor g6795 ( n16559 , n1689 , n26285 );
    or g6796 ( n938 , n29471 , n12668 );
    xnor g6797 ( n21826 , n27453 , n31896 );
    xnor g6798 ( n5349 , n13635 , n8042 );
    and g6799 ( n22378 , n18770 , n22419 );
    and g6800 ( n24039 , n31354 , n22344 );
    xor g6801 ( n1830 , n27098 , n1451 );
    and g6802 ( n834 , n4632 , n747 );
    and g6803 ( n27291 , n30536 , n8975 );
    and g6804 ( n883 , n5145 , n21041 );
    or g6805 ( n4042 , n9120 , n21202 );
    xnor g6806 ( n29801 , n28082 , n17828 );
    xnor g6807 ( n15748 , n8692 , n29457 );
    and g6808 ( n6843 , n29329 , n17009 );
    or g6809 ( n5823 , n24837 , n2801 );
    nor g6810 ( n15799 , n17255 , n26655 );
    or g6811 ( n13068 , n21256 , n12071 );
    or g6812 ( n24211 , n17161 , n2057 );
    and g6813 ( n15393 , n29088 , n5994 );
    xnor g6814 ( n1401 , n2762 , n13764 );
    not g6815 ( n25552 , n25507 );
    xnor g6816 ( n31088 , n25254 , n28441 );
    not g6817 ( n2984 , n17672 );
    or g6818 ( n24188 , n5043 , n30833 );
    not g6819 ( n8610 , n23475 );
    and g6820 ( n16320 , n16013 , n25379 );
    not g6821 ( n24351 , n11270 );
    xnor g6822 ( n30650 , n31970 , n30525 );
    xnor g6823 ( n6647 , n4007 , n31152 );
    or g6824 ( n24051 , n27489 , n10843 );
    nor g6825 ( n27431 , n12668 , n26894 );
    and g6826 ( n22387 , n6441 , n17238 );
    nor g6827 ( n1175 , n19132 , n29746 );
    xnor g6828 ( n20483 , n11954 , n3000 );
    not g6829 ( n7738 , n1521 );
    xnor g6830 ( n19328 , n15532 , n25480 );
    nor g6831 ( n21354 , n11373 , n17981 );
    and g6832 ( n19909 , n16463 , n3737 );
    xnor g6833 ( n24179 , n15919 , n27313 );
    not g6834 ( n25227 , n5949 );
    and g6835 ( n30698 , n17905 , n25977 );
    or g6836 ( n27698 , n14084 , n7679 );
    or g6837 ( n3243 , n5223 , n12278 );
    xnor g6838 ( n27724 , n15638 , n29241 );
    and g6839 ( n29709 , n22428 , n14112 );
    xnor g6840 ( n16654 , n27497 , n25155 );
    and g6841 ( n23814 , n17801 , n10322 );
    nor g6842 ( n13468 , n11313 , n14443 );
    xnor g6843 ( n21680 , n31745 , n27512 );
    xor g6844 ( n27149 , n3135 , n18452 );
    xnor g6845 ( n27356 , n805 , n3347 );
    and g6846 ( n29874 , n6869 , n4236 );
    or g6847 ( n11846 , n5906 , n26438 );
    not g6848 ( n21276 , n19386 );
    nor g6849 ( n21072 , n18650 , n5092 );
    xnor g6850 ( n24272 , n26670 , n14624 );
    not g6851 ( n19888 , n21174 );
    xnor g6852 ( n749 , n28130 , n22194 );
    not g6853 ( n26206 , n29080 );
    not g6854 ( n22563 , n15158 );
    not g6855 ( n31307 , n11964 );
    nor g6856 ( n30816 , n384 , n17352 );
    not g6857 ( n6493 , n18992 );
    and g6858 ( n8880 , n24303 , n4794 );
    nor g6859 ( n20445 , n11247 , n8023 );
    not g6860 ( n18346 , n5806 );
    xnor g6861 ( n893 , n5956 , n29740 );
    nor g6862 ( n26241 , n21606 , n4776 );
    and g6863 ( n29004 , n14886 , n28747 );
    or g6864 ( n10180 , n20155 , n17339 );
    and g6865 ( n19859 , n3222 , n26728 );
    or g6866 ( n25898 , n19475 , n30082 );
    or g6867 ( n11589 , n21169 , n20930 );
    xnor g6868 ( n30424 , n8484 , n26758 );
    nor g6869 ( n7142 , n658 , n21080 );
    xnor g6870 ( n26571 , n20938 , n29886 );
    not g6871 ( n9091 , n30458 );
    or g6872 ( n18137 , n18576 , n12121 );
    nor g6873 ( n20261 , n1036 , n17812 );
    not g6874 ( n18831 , n10519 );
    not g6875 ( n26424 , n10881 );
    xnor g6876 ( n28832 , n26052 , n12055 );
    or g6877 ( n12886 , n12234 , n19019 );
    not g6878 ( n4929 , n17612 );
    or g6879 ( n5402 , n30405 , n25489 );
    or g6880 ( n20134 , n3708 , n7680 );
    not g6881 ( n30617 , n10525 );
    or g6882 ( n29007 , n14191 , n14570 );
    not g6883 ( n11375 , n3259 );
    xnor g6884 ( n14189 , n4012 , n13313 );
    or g6885 ( n29573 , n30699 , n17554 );
    and g6886 ( n12142 , n31375 , n16811 );
    or g6887 ( n22283 , n28687 , n18024 );
    xnor g6888 ( n26447 , n26855 , n7918 );
    not g6889 ( n11238 , n28646 );
    nor g6890 ( n2953 , n6839 , n11469 );
    not g6891 ( n4370 , n30163 );
    not g6892 ( n22927 , n8961 );
    not g6893 ( n31489 , n8869 );
    xnor g6894 ( n15037 , n14449 , n30967 );
    or g6895 ( n21127 , n28734 , n29411 );
    or g6896 ( n25314 , n7834 , n27766 );
    xnor g6897 ( n7770 , n13573 , n14794 );
    not g6898 ( n5665 , n26317 );
    or g6899 ( n17225 , n2595 , n5771 );
    not g6900 ( n27210 , n4311 );
    not g6901 ( n1457 , n26820 );
    or g6902 ( n3834 , n20731 , n12559 );
    not g6903 ( n25808 , n9645 );
    xnor g6904 ( n15083 , n9995 , n12908 );
    not g6905 ( n17184 , n26511 );
    and g6906 ( n3628 , n31461 , n6801 );
    xnor g6907 ( n12026 , n10979 , n29437 );
    nor g6908 ( n11557 , n6745 , n10926 );
    or g6909 ( n2104 , n9586 , n23536 );
    not g6910 ( n29279 , n29993 );
    and g6911 ( n6418 , n860 , n5119 );
    or g6912 ( n67 , n1541 , n30550 );
    xnor g6913 ( n25197 , n19460 , n28638 );
    not g6914 ( n31043 , n15255 );
    and g6915 ( n11690 , n22502 , n2350 );
    and g6916 ( n29550 , n5229 , n25672 );
    nor g6917 ( n7130 , n19590 , n21613 );
    xnor g6918 ( n14064 , n8075 , n27648 );
    not g6919 ( n9574 , n11972 );
    and g6920 ( n10957 , n5933 , n20759 );
    or g6921 ( n3658 , n31510 , n24659 );
    not g6922 ( n25731 , n21212 );
    not g6923 ( n30033 , n20969 );
    and g6924 ( n25285 , n21109 , n9437 );
    or g6925 ( n21845 , n17149 , n29542 );
    nor g6926 ( n28863 , n14589 , n29984 );
    not g6927 ( n18150 , n16776 );
    and g6928 ( n15228 , n26887 , n24429 );
    not g6929 ( n25365 , n30004 );
    and g6930 ( n7333 , n17924 , n27149 );
    xnor g6931 ( n420 , n30482 , n5149 );
    or g6932 ( n17621 , n1878 , n13383 );
    and g6933 ( n10807 , n21398 , n6102 );
    or g6934 ( n27151 , n31420 , n22580 );
    xnor g6935 ( n9036 , n7510 , n20199 );
    and g6936 ( n16960 , n12484 , n20271 );
    xnor g6937 ( n20487 , n2391 , n305 );
    xnor g6938 ( n15379 , n28434 , n1228 );
    or g6939 ( n96 , n24793 , n14357 );
    not g6940 ( n12600 , n8007 );
    not g6941 ( n27131 , n31356 );
    xnor g6942 ( n23485 , n15515 , n12733 );
    or g6943 ( n27611 , n3102 , n6575 );
    xnor g6944 ( n4326 , n2198 , n11470 );
    xnor g6945 ( n2466 , n17311 , n11822 );
    xnor g6946 ( n7999 , n27725 , n25693 );
    xnor g6947 ( n7394 , n29017 , n4607 );
    or g6948 ( n19689 , n1861 , n7344 );
    nor g6949 ( n8912 , n10269 , n20616 );
    xnor g6950 ( n13044 , n23279 , n22159 );
    nor g6951 ( n26667 , n2766 , n29633 );
    or g6952 ( n28071 , n22035 , n773 );
    nor g6953 ( n5146 , n21341 , n18072 );
    xnor g6954 ( n14557 , n32011 , n10034 );
    xnor g6955 ( n27095 , n9416 , n4645 );
    xnor g6956 ( n20183 , n3822 , n11771 );
    or g6957 ( n8079 , n1953 , n27960 );
    and g6958 ( n28162 , n3780 , n15724 );
    or g6959 ( n9678 , n11200 , n26515 );
    or g6960 ( n3017 , n23934 , n18514 );
    or g6961 ( n22758 , n20485 , n28458 );
    or g6962 ( n27905 , n5934 , n7151 );
    and g6963 ( n26550 , n19539 , n27886 );
    not g6964 ( n9176 , n871 );
    xnor g6965 ( n25416 , n30326 , n27534 );
    and g6966 ( n20656 , n17376 , n11581 );
    and g6967 ( n14819 , n11229 , n7660 );
    or g6968 ( n9602 , n28704 , n25847 );
    xnor g6969 ( n31528 , n7844 , n29444 );
    xnor g6970 ( n14012 , n4126 , n5414 );
    and g6971 ( n4473 , n153 , n9409 );
    and g6972 ( n16144 , n7996 , n1640 );
    not g6973 ( n20793 , n15363 );
    or g6974 ( n11882 , n14154 , n26938 );
    or g6975 ( n1080 , n15397 , n5834 );
    and g6976 ( n18699 , n11534 , n15263 );
    not g6977 ( n2005 , n14087 );
    xnor g6978 ( n2615 , n3824 , n31255 );
    or g6979 ( n23729 , n10936 , n15446 );
    or g6980 ( n9041 , n6586 , n24836 );
    xnor g6981 ( n20074 , n4260 , n9427 );
    not g6982 ( n929 , n30174 );
    xnor g6983 ( n974 , n10988 , n30564 );
    xnor g6984 ( n24161 , n13774 , n7910 );
    and g6985 ( n29012 , n5393 , n6158 );
    not g6986 ( n30955 , n13677 );
    or g6987 ( n13873 , n16568 , n5932 );
    not g6988 ( n29039 , n8988 );
    not g6989 ( n7466 , n24138 );
    xnor g6990 ( n28287 , n18389 , n4213 );
    or g6991 ( n2796 , n17788 , n16025 );
    xor g6992 ( n15232 , n25708 , n10801 );
    and g6993 ( n25455 , n15175 , n27921 );
    not g6994 ( n24828 , n23557 );
    not g6995 ( n28947 , n24243 );
    and g6996 ( n10336 , n19894 , n18484 );
    not g6997 ( n2256 , n3795 );
    or g6998 ( n16206 , n16729 , n26496 );
    xnor g6999 ( n3221 , n31248 , n11262 );
    or g7000 ( n18998 , n15941 , n23942 );
    xnor g7001 ( n17536 , n31412 , n12261 );
    not g7002 ( n31928 , n26298 );
    nor g7003 ( n30220 , n27805 , n6804 );
    nor g7004 ( n10063 , n8388 , n9806 );
    xnor g7005 ( n20507 , n5382 , n26619 );
    and g7006 ( n18359 , n13565 , n28349 );
    xnor g7007 ( n30378 , n3659 , n11985 );
    not g7008 ( n16357 , n8834 );
    and g7009 ( n30666 , n20229 , n14898 );
    xnor g7010 ( n329 , n28202 , n16120 );
    not g7011 ( n14488 , n7465 );
    xor g7012 ( n4951 , n23948 , n24988 );
    and g7013 ( n26455 , n13553 , n22295 );
    not g7014 ( n22737 , n24165 );
    not g7015 ( n19575 , n15376 );
    not g7016 ( n28127 , n2675 );
    or g7017 ( n30463 , n5061 , n8687 );
    buf g7018 ( n11648 , n31000 );
    xnor g7019 ( n28225 , n5352 , n26260 );
    and g7020 ( n1244 , n22092 , n24302 );
    and g7021 ( n6159 , n1249 , n7832 );
    xnor g7022 ( n5288 , n6032 , n16755 );
    not g7023 ( n23607 , n16608 );
    not g7024 ( n1476 , n17572 );
    not g7025 ( n22203 , n17851 );
    and g7026 ( n18854 , n17050 , n15011 );
    and g7027 ( n6050 , n4722 , n14967 );
    xnor g7028 ( n3579 , n17963 , n11265 );
    and g7029 ( n6052 , n2644 , n1219 );
    xnor g7030 ( n9783 , n28846 , n23154 );
    nor g7031 ( n7647 , n16790 , n31781 );
    or g7032 ( n8594 , n7390 , n29190 );
    not g7033 ( n11037 , n9445 );
    not g7034 ( n23456 , n21793 );
    not g7035 ( n31492 , n5313 );
    xnor g7036 ( n29611 , n1291 , n4936 );
    not g7037 ( n22631 , n16516 );
    or g7038 ( n20297 , n27975 , n9638 );
    nor g7039 ( n11684 , n13733 , n16256 );
    nor g7040 ( n6935 , n13517 , n10794 );
    or g7041 ( n6231 , n22241 , n6095 );
    nor g7042 ( n7350 , n4847 , n12207 );
    nor g7043 ( n30342 , n13833 , n18506 );
    or g7044 ( n25729 , n27857 , n29531 );
    or g7045 ( n4772 , n4836 , n13708 );
    or g7046 ( n26829 , n1208 , n24328 );
    or g7047 ( n8958 , n14001 , n29288 );
    not g7048 ( n11319 , n14201 );
    nor g7049 ( n29203 , n15758 , n13833 );
    xnor g7050 ( n30177 , n21771 , n26996 );
    xnor g7051 ( n21281 , n31423 , n28738 );
    nor g7052 ( n10577 , n10665 , n18454 );
    not g7053 ( n8918 , n23720 );
    xnor g7054 ( n11995 , n5348 , n24738 );
    xnor g7055 ( n16275 , n9713 , n24617 );
    or g7056 ( n20651 , n7923 , n8729 );
    or g7057 ( n11659 , n21638 , n10223 );
    or g7058 ( n30430 , n16706 , n28212 );
    not g7059 ( n2127 , n9162 );
    xnor g7060 ( n7439 , n16004 , n5004 );
    and g7061 ( n18779 , n5410 , n16462 );
    not g7062 ( n8602 , n3636 );
    and g7063 ( n23265 , n25151 , n7961 );
    not g7064 ( n29063 , n25994 );
    not g7065 ( n6166 , n15232 );
    xnor g7066 ( n31320 , n25584 , n707 );
    and g7067 ( n4497 , n5005 , n13731 );
    or g7068 ( n4082 , n23052 , n20622 );
    or g7069 ( n7449 , n12697 , n24560 );
    xnor g7070 ( n30181 , n1132 , n840 );
    xnor g7071 ( n27274 , n21075 , n16452 );
    xnor g7072 ( n29996 , n25706 , n14741 );
    or g7073 ( n27130 , n14315 , n14561 );
    not g7074 ( n21070 , n26464 );
    and g7075 ( n11014 , n16075 , n15588 );
    xnor g7076 ( n4023 , n29877 , n2004 );
    not g7077 ( n16300 , n23643 );
    xnor g7078 ( n25689 , n31364 , n6304 );
    and g7079 ( n15117 , n27548 , n10303 );
    and g7080 ( n22060 , n14743 , n7998 );
    not g7081 ( n29578 , n14024 );
    not g7082 ( n5985 , n23521 );
    xor g7083 ( n22357 , n26854 , n2681 );
    xnor g7084 ( n18839 , n30975 , n20379 );
    or g7085 ( n10816 , n21599 , n21360 );
    or g7086 ( n8825 , n23040 , n8834 );
    or g7087 ( n12984 , n13052 , n24994 );
    not g7088 ( n5441 , n29444 );
    not g7089 ( n8232 , n6003 );
    or g7090 ( n13139 , n12632 , n30388 );
    or g7091 ( n27809 , n6459 , n31392 );
    xnor g7092 ( n31617 , n18180 , n643 );
    or g7093 ( n6463 , n14954 , n12396 );
    or g7094 ( n26883 , n8107 , n29456 );
    not g7095 ( n21579 , n22450 );
    or g7096 ( n28380 , n5204 , n11865 );
    or g7097 ( n23091 , n22226 , n24949 );
    xnor g7098 ( n7789 , n14856 , n4509 );
    xnor g7099 ( n15265 , n20632 , n561 );
    and g7100 ( n17012 , n31899 , n4689 );
    and g7101 ( n22110 , n24438 , n6235 );
    and g7102 ( n10858 , n25054 , n992 );
    not g7103 ( n24964 , n26859 );
    or g7104 ( n8230 , n1635 , n28260 );
    and g7105 ( n23864 , n23688 , n2101 );
    or g7106 ( n16973 , n13295 , n4701 );
    not g7107 ( n6087 , n4210 );
    not g7108 ( n10380 , n29259 );
    xnor g7109 ( n13559 , n9378 , n3930 );
    or g7110 ( n14886 , n12167 , n23150 );
    not g7111 ( n16642 , n9490 );
    xor g7112 ( n29963 , n15866 , n8091 );
    or g7113 ( n25815 , n19061 , n14919 );
    or g7114 ( n12436 , n355 , n15180 );
    not g7115 ( n14808 , n9551 );
    xnor g7116 ( n28395 , n3166 , n4847 );
    not g7117 ( n21019 , n22917 );
    not g7118 ( n26239 , n21377 );
    and g7119 ( n23637 , n2016 , n10748 );
    or g7120 ( n756 , n24043 , n28702 );
    and g7121 ( n19370 , n23461 , n7669 );
    xnor g7122 ( n8320 , n1762 , n5965 );
    and g7123 ( n24216 , n23346 , n24323 );
    not g7124 ( n23491 , n5560 );
    and g7125 ( n8409 , n13620 , n22593 );
    xnor g7126 ( n30975 , n17377 , n1792 );
    and g7127 ( n9617 , n28566 , n28607 );
    and g7128 ( n20207 , n21744 , n12864 );
    or g7129 ( n27393 , n31916 , n14831 );
    xnor g7130 ( n2287 , n7020 , n24564 );
    not g7131 ( n2688 , n28141 );
    or g7132 ( n31383 , n1762 , n12716 );
    not g7133 ( n25864 , n26786 );
    xnor g7134 ( n25741 , n7240 , n18734 );
    xnor g7135 ( n1808 , n13561 , n30431 );
    xnor g7136 ( n15785 , n20580 , n15112 );
    not g7137 ( n13949 , n9655 );
    xnor g7138 ( n4020 , n11692 , n20736 );
    not g7139 ( n493 , n9760 );
    not g7140 ( n9609 , n1260 );
    nor g7141 ( n25817 , n10477 , n683 );
    xnor g7142 ( n7059 , n1067 , n5561 );
    xnor g7143 ( n16917 , n19531 , n21340 );
    nor g7144 ( n29869 , n26625 , n21560 );
    not g7145 ( n2687 , n17189 );
    not g7146 ( n12784 , n2271 );
    xnor g7147 ( n29382 , n10575 , n4593 );
    not g7148 ( n6359 , n9706 );
    xnor g7149 ( n20560 , n23606 , n30753 );
    not g7150 ( n28332 , n1480 );
    not g7151 ( n29343 , n8173 );
    and g7152 ( n3784 , n5167 , n1001 );
    or g7153 ( n6227 , n27336 , n28379 );
    or g7154 ( n13469 , n13023 , n22998 );
    and g7155 ( n6911 , n26544 , n1980 );
    xnor g7156 ( n620 , n2374 , n15286 );
    xnor g7157 ( n12799 , n19615 , n12210 );
    nor g7158 ( n15270 , n2301 , n30948 );
    not g7159 ( n2437 , n29710 );
    xnor g7160 ( n16240 , n22842 , n9691 );
    nor g7161 ( n4649 , n7098 , n7137 );
    xnor g7162 ( n10242 , n3335 , n16061 );
    xnor g7163 ( n27553 , n19960 , n31306 );
    or g7164 ( n14050 , n24474 , n1468 );
    xnor g7165 ( n10917 , n18489 , n1285 );
    or g7166 ( n30138 , n27343 , n2232 );
    or g7167 ( n28385 , n19845 , n15539 );
    xnor g7168 ( n23406 , n207 , n25380 );
    xnor g7169 ( n4949 , n30891 , n27978 );
    and g7170 ( n6495 , n9006 , n7302 );
    xnor g7171 ( n14109 , n8249 , n22852 );
    or g7172 ( n18814 , n22172 , n17834 );
    buf g7173 ( n3269 , n4952 );
    or g7174 ( n26782 , n30221 , n6749 );
    and g7175 ( n14169 , n18046 , n26986 );
    nor g7176 ( n20831 , n661 , n22275 );
    xnor g7177 ( n20889 , n8577 , n22512 );
    and g7178 ( n28309 , n30613 , n28263 );
    or g7179 ( n19667 , n8693 , n13655 );
    nor g7180 ( n20064 , n10013 , n32028 );
    not g7181 ( n7552 , n12713 );
    nor g7182 ( n22939 , n6534 , n21589 );
    nor g7183 ( n20027 , n7720 , n9190 );
    xnor g7184 ( n1708 , n3438 , n24876 );
    xor g7185 ( n10793 , n8506 , n18001 );
    or g7186 ( n6290 , n9744 , n22841 );
    not g7187 ( n27213 , n6701 );
    not g7188 ( n11911 , n8492 );
    not g7189 ( n5305 , n17617 );
    not g7190 ( n18208 , n31232 );
    and g7191 ( n6408 , n2327 , n217 );
    not g7192 ( n25997 , n12668 );
    or g7193 ( n27263 , n26512 , n3034 );
    or g7194 ( n19047 , n4371 , n3083 );
    and g7195 ( n12579 , n25207 , n23836 );
    nor g7196 ( n24488 , n12979 , n31369 );
    xnor g7197 ( n389 , n23561 , n22233 );
    or g7198 ( n3741 , n8641 , n19705 );
    not g7199 ( n4747 , n26743 );
    xnor g7200 ( n16619 , n20814 , n9361 );
    not g7201 ( n1787 , n28111 );
    not g7202 ( n26331 , n1275 );
    and g7203 ( n19613 , n27607 , n26857 );
    not g7204 ( n21882 , n22974 );
    or g7205 ( n16501 , n7228 , n10441 );
    and g7206 ( n26305 , n4078 , n21763 );
    and g7207 ( n30038 , n16928 , n23703 );
    not g7208 ( n13375 , n20987 );
    buf g7209 ( n25798 , n10229 );
    not g7210 ( n7456 , n14518 );
    xnor g7211 ( n5883 , n24265 , n27597 );
    or g7212 ( n2907 , n12613 , n29330 );
    xnor g7213 ( n18958 , n19892 , n9744 );
    xnor g7214 ( n26525 , n12389 , n28395 );
    not g7215 ( n15726 , n19817 );
    not g7216 ( n33 , n1177 );
    and g7217 ( n3796 , n30261 , n1659 );
    not g7218 ( n9626 , n19765 );
    xnor g7219 ( n5633 , n12357 , n30337 );
    xnor g7220 ( n28965 , n28576 , n23485 );
    not g7221 ( n13352 , n2638 );
    or g7222 ( n22950 , n8794 , n9315 );
    or g7223 ( n13775 , n27476 , n9770 );
    and g7224 ( n8447 , n240 , n28264 );
    not g7225 ( n23064 , n15941 );
    or g7226 ( n31871 , n19592 , n28683 );
    and g7227 ( n25824 , n11311 , n9991 );
    and g7228 ( n22351 , n12594 , n1078 );
    xnor g7229 ( n14105 , n10970 , n18544 );
    xnor g7230 ( n17460 , n29551 , n19011 );
    or g7231 ( n24809 , n23014 , n18466 );
    and g7232 ( n10057 , n8569 , n6765 );
    or g7233 ( n26394 , n29378 , n854 );
    and g7234 ( n30333 , n13428 , n9937 );
    xnor g7235 ( n9280 , n22156 , n13342 );
    or g7236 ( n9436 , n14992 , n41 );
    xnor g7237 ( n8493 , n30463 , n8487 );
    xnor g7238 ( n11907 , n6576 , n27427 );
    not g7239 ( n22687 , n7409 );
    xnor g7240 ( n26001 , n26766 , n3880 );
    xnor g7241 ( n8784 , n6545 , n20060 );
    xnor g7242 ( n13786 , n30465 , n27196 );
    not g7243 ( n10108 , n1304 );
    and g7244 ( n17982 , n31697 , n14957 );
    xnor g7245 ( n6027 , n19483 , n21968 );
    xnor g7246 ( n27472 , n30261 , n26817 );
    or g7247 ( n22436 , n3450 , n10555 );
    xnor g7248 ( n27806 , n29933 , n11361 );
    nor g7249 ( n21592 , n23679 , n18848 );
    xnor g7250 ( n29630 , n27829 , n1039 );
    and g7251 ( n25772 , n9331 , n22478 );
    xnor g7252 ( n7080 , n22107 , n11801 );
    not g7253 ( n7039 , n30872 );
    nor g7254 ( n12062 , n9639 , n9579 );
    not g7255 ( n12720 , n16659 );
    nor g7256 ( n15894 , n6249 , n31170 );
    xnor g7257 ( n30768 , n24423 , n19211 );
    and g7258 ( n19836 , n12512 , n3748 );
    nor g7259 ( n20983 , n21258 , n10414 );
    and g7260 ( n18454 , n841 , n25696 );
    not g7261 ( n12412 , n18852 );
    or g7262 ( n7167 , n9844 , n10324 );
    or g7263 ( n26152 , n29198 , n29772 );
    or g7264 ( n17668 , n5758 , n3388 );
    and g7265 ( n31478 , n6022 , n19115 );
    or g7266 ( n23768 , n19929 , n14982 );
    not g7267 ( n7 , n11543 );
    xnor g7268 ( n14667 , n27074 , n24958 );
    not g7269 ( n5314 , n5525 );
    xnor g7270 ( n1109 , n26965 , n2375 );
    xnor g7271 ( n2784 , n13145 , n9935 );
    not g7272 ( n14391 , n2231 );
    nor g7273 ( n8490 , n26052 , n7471 );
    xnor g7274 ( n2417 , n16347 , n18002 );
    not g7275 ( n9994 , n8936 );
    xnor g7276 ( n31376 , n6464 , n4468 );
    not g7277 ( n24442 , n16922 );
    nor g7278 ( n14153 , n6172 , n25818 );
    or g7279 ( n31551 , n7566 , n5336 );
    not g7280 ( n25792 , n8545 );
    xnor g7281 ( n15144 , n844 , n20889 );
    and g7282 ( n12389 , n17049 , n18665 );
    nor g7283 ( n12568 , n14926 , n2845 );
    xor g7284 ( n812 , n9660 , n30936 );
    or g7285 ( n11664 , n3022 , n15094 );
    nor g7286 ( n15237 , n28781 , n29891 );
    xnor g7287 ( n29905 , n4648 , n833 );
    not g7288 ( n3210 , n1935 );
    or g7289 ( n12291 , n25098 , n4589 );
    or g7290 ( n7388 , n23647 , n25627 );
    xnor g7291 ( n4165 , n6162 , n19536 );
    and g7292 ( n20992 , n25944 , n9249 );
    nor g7293 ( n31293 , n29578 , n14380 );
    and g7294 ( n27520 , n20110 , n16340 );
    not g7295 ( n5047 , n25398 );
    nor g7296 ( n8416 , n31514 , n17024 );
    and g7297 ( n20481 , n7497 , n8422 );
    xnor g7298 ( n19986 , n21115 , n14906 );
    xnor g7299 ( n31455 , n16144 , n1712 );
    not g7300 ( n31809 , n10880 );
    and g7301 ( n4544 , n8743 , n13956 );
    or g7302 ( n3556 , n23677 , n24356 );
    or g7303 ( n16878 , n3479 , n70 );
    not g7304 ( n9351 , n25169 );
    or g7305 ( n23753 , n30102 , n22841 );
    not g7306 ( n11339 , n8760 );
    not g7307 ( n3743 , n16593 );
    or g7308 ( n15461 , n16509 , n20936 );
    xnor g7309 ( n18116 , n27609 , n3837 );
    xnor g7310 ( n17048 , n9396 , n31094 );
    xnor g7311 ( n726 , n18825 , n4054 );
    not g7312 ( n601 , n29678 );
    and g7313 ( n19213 , n29018 , n19438 );
    not g7314 ( n17860 , n11692 );
    and g7315 ( n17337 , n14202 , n4956 );
    xnor g7316 ( n8197 , n3822 , n7414 );
    not g7317 ( n5710 , n19107 );
    xnor g7318 ( n6779 , n25204 , n20740 );
    xnor g7319 ( n24431 , n1509 , n412 );
    or g7320 ( n25811 , n29569 , n1871 );
    xnor g7321 ( n31623 , n3879 , n28466 );
    xnor g7322 ( n22118 , n28553 , n18793 );
    and g7323 ( n5111 , n27165 , n20624 );
    or g7324 ( n19028 , n18248 , n14472 );
    xnor g7325 ( n3347 , n16412 , n2597 );
    and g7326 ( n19016 , n10182 , n14687 );
    xnor g7327 ( n20763 , n31049 , n22244 );
    not g7328 ( n4610 , n13749 );
    not g7329 ( n22172 , n30522 );
    not g7330 ( n18104 , n27301 );
    not g7331 ( n23947 , n5411 );
    not g7332 ( n26743 , n23485 );
    not g7333 ( n11244 , n7692 );
    xnor g7334 ( n14246 , n787 , n10477 );
    xor g7335 ( n515 , n383 , n11051 );
    or g7336 ( n22502 , n16390 , n10679 );
    and g7337 ( n21619 , n29863 , n21123 );
    xnor g7338 ( n7796 , n5972 , n11592 );
    xnor g7339 ( n6454 , n19471 , n16603 );
    xnor g7340 ( n18624 , n6554 , n14098 );
    or g7341 ( n13742 , n26933 , n30693 );
    xor g7342 ( n31277 , n5103 , n8567 );
    not g7343 ( n15635 , n17338 );
    not g7344 ( n5902 , n8669 );
    not g7345 ( n10636 , n7254 );
    xnor g7346 ( n30907 , n30156 , n19214 );
    not g7347 ( n18524 , n18537 );
    xnor g7348 ( n21801 , n26857 , n5052 );
    or g7349 ( n15498 , n27385 , n25565 );
    not g7350 ( n29305 , n8852 );
    or g7351 ( n18567 , n1004 , n23554 );
    xnor g7352 ( n30794 , n8624 , n30908 );
    nor g7353 ( n5444 , n11771 , n16689 );
    or g7354 ( n29179 , n28621 , n11740 );
    not g7355 ( n3064 , n7470 );
    and g7356 ( n11203 , n19243 , n19561 );
    or g7357 ( n1259 , n4877 , n29148 );
    nor g7358 ( n11776 , n9591 , n9137 );
    or g7359 ( n13341 , n13960 , n8695 );
    xnor g7360 ( n22649 , n5115 , n12201 );
    and g7361 ( n2890 , n10766 , n26111 );
    not g7362 ( n4135 , n15680 );
    and g7363 ( n18310 , n16792 , n18392 );
    and g7364 ( n3097 , n15104 , n11762 );
    xnor g7365 ( n9980 , n25878 , n1679 );
    nor g7366 ( n17168 , n24118 , n2798 );
    or g7367 ( n9958 , n28065 , n2439 );
    not g7368 ( n9879 , n2292 );
    nor g7369 ( n27025 , n19378 , n30504 );
    not g7370 ( n27827 , n6965 );
    not g7371 ( n16575 , n22340 );
    not g7372 ( n13797 , n30444 );
    and g7373 ( n4081 , n14685 , n3964 );
    or g7374 ( n8651 , n8861 , n24843 );
    xnor g7375 ( n21717 , n10679 , n31948 );
    xnor g7376 ( n21706 , n27800 , n5650 );
    xnor g7377 ( n12530 , n5748 , n13012 );
    or g7378 ( n25191 , n14747 , n11377 );
    nor g7379 ( n1257 , n28270 , n7090 );
    or g7380 ( n28997 , n851 , n8601 );
    not g7381 ( n18149 , n21032 );
    and g7382 ( n23180 , n14347 , n9454 );
    xor g7383 ( n25284 , n8283 , n758 );
    not g7384 ( n25252 , n9530 );
    xnor g7385 ( n951 , n14428 , n22029 );
    or g7386 ( n16662 , n2508 , n8776 );
    and g7387 ( n17456 , n31236 , n23286 );
    buf g7388 ( n28445 , n8563 );
    and g7389 ( n440 , n3996 , n16856 );
    not g7390 ( n20878 , n30198 );
    or g7391 ( n22102 , n3837 , n17847 );
    buf g7392 ( n31918 , n10398 );
    or g7393 ( n14762 , n3042 , n7375 );
    or g7394 ( n22786 , n14865 , n15205 );
    nor g7395 ( n20195 , n19384 , n11002 );
    xnor g7396 ( n15901 , n15818 , n20210 );
    and g7397 ( n10518 , n16817 , n11828 );
    nor g7398 ( n23075 , n5401 , n17931 );
    xor g7399 ( n17762 , n9169 , n6803 );
    not g7400 ( n11998 , n1669 );
    not g7401 ( n17904 , n27520 );
    nor g7402 ( n984 , n23366 , n19859 );
    xnor g7403 ( n31643 , n30349 , n10269 );
    not g7404 ( n20149 , n13092 );
    not g7405 ( n4939 , n22352 );
    not g7406 ( n9056 , n30681 );
    xnor g7407 ( n8418 , n29653 , n6179 );
    not g7408 ( n15161 , n29559 );
    not g7409 ( n30254 , n8321 );
    not g7410 ( n20856 , n24032 );
    and g7411 ( n22583 , n23147 , n20138 );
    not g7412 ( n31023 , n23311 );
    not g7413 ( n14901 , n22521 );
    not g7414 ( n2289 , n18671 );
    and g7415 ( n9271 , n17264 , n19418 );
    or g7416 ( n27050 , n8469 , n28992 );
    not g7417 ( n7050 , n28580 );
    and g7418 ( n13668 , n24476 , n26078 );
    or g7419 ( n7952 , n30558 , n978 );
    xnor g7420 ( n20342 , n28829 , n5022 );
    xnor g7421 ( n3416 , n30890 , n8986 );
    and g7422 ( n17406 , n18788 , n4498 );
    not g7423 ( n23559 , n29663 );
    and g7424 ( n28596 , n20694 , n3031 );
    xnor g7425 ( n18947 , n6667 , n23561 );
    buf g7426 ( n19892 , n5275 );
    or g7427 ( n25662 , n2560 , n1642 );
    xnor g7428 ( n30814 , n20453 , n30769 );
    or g7429 ( n7480 , n9326 , n13119 );
    not g7430 ( n23949 , n16387 );
    xnor g7431 ( n28464 , n22197 , n11905 );
    xnor g7432 ( n14454 , n17286 , n12006 );
    nor g7433 ( n17106 , n10158 , n18503 );
    or g7434 ( n24796 , n15191 , n5847 );
    xnor g7435 ( n1365 , n485 , n27243 );
    or g7436 ( n28307 , n29169 , n13892 );
    and g7437 ( n29942 , n14436 , n21351 );
    xnor g7438 ( n15298 , n1456 , n21850 );
    xnor g7439 ( n18725 , n14829 , n9010 );
    and g7440 ( n6769 , n24502 , n6001 );
    xnor g7441 ( n25219 , n11699 , n2336 );
    not g7442 ( n12041 , n23498 );
    or g7443 ( n17502 , n5959 , n17978 );
    not g7444 ( n14738 , n9266 );
    not g7445 ( n20192 , n32001 );
    not g7446 ( n9886 , n31857 );
    or g7447 ( n647 , n5665 , n20705 );
    nor g7448 ( n6657 , n12399 , n7473 );
    not g7449 ( n22251 , n8969 );
    not g7450 ( n1696 , n30505 );
    buf g7451 ( n30227 , n17110 );
    xnor g7452 ( n13602 , n4354 , n27325 );
    or g7453 ( n18663 , n15558 , n9435 );
    xnor g7454 ( n7993 , n20412 , n11360 );
    and g7455 ( n16962 , n31752 , n27927 );
    and g7456 ( n14339 , n11369 , n558 );
    or g7457 ( n7135 , n11708 , n15662 );
    or g7458 ( n4290 , n29029 , n9514 );
    or g7459 ( n5993 , n21265 , n27012 );
    xnor g7460 ( n10471 , n3255 , n12154 );
    not g7461 ( n16002 , n5789 );
    not g7462 ( n2679 , n21508 );
    nor g7463 ( n23887 , n27848 , n25176 );
    xnor g7464 ( n4881 , n6086 , n2558 );
    not g7465 ( n24459 , n22233 );
    or g7466 ( n3543 , n23695 , n20281 );
    xnor g7467 ( n16963 , n23371 , n5725 );
    xnor g7468 ( n11155 , n8461 , n5454 );
    or g7469 ( n29675 , n8184 , n29498 );
    nor g7470 ( n13947 , n14954 , n17611 );
    xnor g7471 ( n31482 , n30908 , n20236 );
    and g7472 ( n873 , n28959 , n10587 );
    or g7473 ( n15003 , n17871 , n9119 );
    not g7474 ( n8089 , n8054 );
    and g7475 ( n21324 , n20471 , n25773 );
    or g7476 ( n31045 , n9456 , n7887 );
    and g7477 ( n1656 , n26017 , n24951 );
    xnor g7478 ( n19631 , n333 , n29051 );
    or g7479 ( n18176 , n6139 , n5825 );
    xnor g7480 ( n23614 , n6781 , n29276 );
    or g7481 ( n8458 , n24459 , n9538 );
    or g7482 ( n2974 , n12700 , n1296 );
    and g7483 ( n3736 , n8233 , n26640 );
    or g7484 ( n4076 , n17169 , n14819 );
    and g7485 ( n31159 , n8692 , n10180 );
    or g7486 ( n18459 , n12840 , n23316 );
    or g7487 ( n1793 , n15558 , n24464 );
    not g7488 ( n222 , n25066 );
    or g7489 ( n26498 , n25860 , n14082 );
    xnor g7490 ( n11654 , n3765 , n238 );
    or g7491 ( n28865 , n21027 , n12852 );
    and g7492 ( n9542 , n5958 , n9997 );
    and g7493 ( n14650 , n15546 , n19321 );
    or g7494 ( n23139 , n28191 , n16974 );
    nor g7495 ( n13224 , n8815 , n18668 );
    or g7496 ( n17629 , n4584 , n25931 );
    or g7497 ( n24629 , n3254 , n16218 );
    or g7498 ( n10725 , n5022 , n30323 );
    nor g7499 ( n7512 , n16075 , n30201 );
    nor g7500 ( n27598 , n144 , n17107 );
    nor g7501 ( n8259 , n1742 , n19317 );
    xnor g7502 ( n19316 , n13137 , n27805 );
    not g7503 ( n21537 , n5598 );
    not g7504 ( n2646 , n17291 );
    xnor g7505 ( n21655 , n17075 , n29317 );
    and g7506 ( n18934 , n9363 , n13245 );
    or g7507 ( n16644 , n18899 , n4643 );
    xnor g7508 ( n29661 , n18834 , n24127 );
    xnor g7509 ( n3921 , n19405 , n17499 );
    or g7510 ( n17140 , n14631 , n19086 );
    or g7511 ( n16985 , n11005 , n6539 );
    nor g7512 ( n1723 , n29153 , n18808 );
    xnor g7513 ( n13912 , n5923 , n7732 );
    or g7514 ( n20048 , n16261 , n10777 );
    or g7515 ( n5919 , n8449 , n10241 );
    xnor g7516 ( n14107 , n7434 , n22512 );
    or g7517 ( n6501 , n11462 , n14147 );
    xnor g7518 ( n5211 , n19886 , n817 );
    xnor g7519 ( n31456 , n12477 , n15845 );
    not g7520 ( n15662 , n6590 );
    and g7521 ( n18736 , n9594 , n7203 );
    xnor g7522 ( n9115 , n26144 , n6178 );
    xnor g7523 ( n22470 , n22518 , n9173 );
    nor g7524 ( n21937 , n7425 , n15776 );
    or g7525 ( n24701 , n17279 , n1893 );
    nor g7526 ( n22247 , n2435 , n31256 );
    or g7527 ( n21483 , n20539 , n31717 );
    not g7528 ( n14742 , n22114 );
    xnor g7529 ( n31924 , n10619 , n14324 );
    not g7530 ( n17235 , n12683 );
    nor g7531 ( n10580 , n14828 , n20625 );
    not g7532 ( n24639 , n29902 );
    and g7533 ( n12657 , n322 , n30687 );
    xnor g7534 ( n2913 , n8049 , n18507 );
    nor g7535 ( n30905 , n17851 , n2263 );
    not g7536 ( n29083 , n10870 );
    not g7537 ( n8390 , n20141 );
    not g7538 ( n5380 , n24766 );
    not g7539 ( n21116 , n20660 );
    not g7540 ( n26468 , n26923 );
    not g7541 ( n14842 , n12422 );
    not g7542 ( n6927 , n4777 );
    or g7543 ( n13182 , n895 , n4363 );
    and g7544 ( n23717 , n10950 , n25166 );
    xnor g7545 ( n30474 , n14708 , n16106 );
    not g7546 ( n31535 , n14105 );
    not g7547 ( n19593 , n9391 );
    or g7548 ( n21652 , n7180 , n27121 );
    not g7549 ( n10557 , n3461 );
    xnor g7550 ( n23208 , n27602 , n23828 );
    and g7551 ( n22998 , n22524 , n23416 );
    and g7552 ( n11382 , n5544 , n30623 );
    or g7553 ( n25268 , n1656 , n14058 );
    nor g7554 ( n14526 , n22845 , n1670 );
    or g7555 ( n6252 , n19864 , n8522 );
    not g7556 ( n3915 , n31419 );
    not g7557 ( n16092 , n20202 );
    or g7558 ( n9102 , n7707 , n12706 );
    not g7559 ( n28576 , n10197 );
    or g7560 ( n16713 , n6803 , n9169 );
    and g7561 ( n7684 , n5946 , n13687 );
    xnor g7562 ( n18282 , n10027 , n18924 );
    or g7563 ( n5000 , n15466 , n29869 );
    nor g7564 ( n26245 , n18507 , n11340 );
    and g7565 ( n3398 , n13001 , n4980 );
    or g7566 ( n15650 , n16082 , n6843 );
    not g7567 ( n2368 , n24570 );
    or g7568 ( n30696 , n12494 , n11167 );
    nor g7569 ( n18899 , n20043 , n7535 );
    and g7570 ( n29544 , n30652 , n29193 );
    not g7571 ( n18418 , n29305 );
    nor g7572 ( n28874 , n28006 , n5149 );
    xor g7573 ( n22907 , n19909 , n19562 );
    or g7574 ( n21650 , n27504 , n4382 );
    and g7575 ( n10110 , n4390 , n6799 );
    and g7576 ( n29848 , n31220 , n14972 );
    not g7577 ( n14366 , n5270 );
    and g7578 ( n16335 , n25685 , n1160 );
    not g7579 ( n26312 , n30165 );
    xor g7580 ( n7812 , n31175 , n31213 );
    or g7581 ( n2838 , n10334 , n669 );
    xnor g7582 ( n807 , n29800 , n28533 );
    not g7583 ( n18800 , n6780 );
    not g7584 ( n26069 , n12593 );
    not g7585 ( n15577 , n4446 );
    or g7586 ( n14142 , n28231 , n15970 );
    xnor g7587 ( n31104 , n28689 , n11422 );
    or g7588 ( n27114 , n31326 , n3902 );
    nor g7589 ( n14689 , n27804 , n12117 );
    nor g7590 ( n30836 , n23115 , n16075 );
    not g7591 ( n13212 , n1940 );
    nor g7592 ( n3840 , n5358 , n30686 );
    not g7593 ( n15452 , n4130 );
    xor g7594 ( n24210 , n28778 , n8447 );
    and g7595 ( n8598 , n13353 , n14540 );
    not g7596 ( n5268 , n6404 );
    and g7597 ( n13641 , n11699 , n30537 );
    xnor g7598 ( n8782 , n25191 , n30026 );
    not g7599 ( n5901 , n3471 );
    nor g7600 ( n242 , n23153 , n24063 );
    not g7601 ( n23109 , n27994 );
    not g7602 ( n20754 , n19422 );
    or g7603 ( n1310 , n29993 , n1587 );
    nor g7604 ( n12552 , n7240 , n12405 );
    not g7605 ( n11472 , n31652 );
    xnor g7606 ( n28738 , n11157 , n22549 );
    xnor g7607 ( n23720 , n1075 , n10836 );
    not g7608 ( n28370 , n24916 );
    and g7609 ( n3215 , n23625 , n14326 );
    not g7610 ( n8107 , n5350 );
    or g7611 ( n11449 , n18955 , n6072 );
    and g7612 ( n11088 , n13315 , n8956 );
    not g7613 ( n20626 , n29274 );
    not g7614 ( n6240 , n22561 );
    and g7615 ( n30319 , n3517 , n19165 );
    or g7616 ( n19595 , n18253 , n23119 );
    not g7617 ( n5328 , n17038 );
    or g7618 ( n31724 , n15053 , n14314 );
    not g7619 ( n25709 , n21723 );
    xnor g7620 ( n24093 , n9940 , n3388 );
    not g7621 ( n5816 , n6160 );
    or g7622 ( n11966 , n28879 , n13730 );
    xor g7623 ( n27390 , n17198 , n5846 );
    or g7624 ( n19050 , n7559 , n18902 );
    or g7625 ( n25406 , n27906 , n4451 );
    not g7626 ( n25 , n2666 );
    nor g7627 ( n1854 , n3372 , n22268 );
    not g7628 ( n3971 , n3963 );
    not g7629 ( n19946 , n14363 );
    not g7630 ( n28686 , n13514 );
    not g7631 ( n12675 , n26792 );
    nor g7632 ( n9646 , n5190 , n1284 );
    nor g7633 ( n14675 , n23561 , n20663 );
    not g7634 ( n4045 , n23419 );
    or g7635 ( n414 , n1600 , n24630 );
    not g7636 ( n10550 , n14484 );
    xnor g7637 ( n31375 , n3344 , n26227 );
    not g7638 ( n30420 , n24256 );
    and g7639 ( n31501 , n14483 , n3922 );
    buf g7640 ( n17771 , n21643 );
    and g7641 ( n18774 , n9347 , n4585 );
    not g7642 ( n12825 , n18425 );
    and g7643 ( n6710 , n2380 , n20745 );
    not g7644 ( n3412 , n3858 );
    not g7645 ( n1094 , n30040 );
    xnor g7646 ( n31042 , n5995 , n26561 );
    and g7647 ( n16416 , n31172 , n560 );
    nor g7648 ( n17259 , n5288 , n14280 );
    and g7649 ( n4546 , n313 , n28255 );
    or g7650 ( n4746 , n26544 , n19315 );
    or g7651 ( n7856 , n688 , n22952 );
    not g7652 ( n4524 , n3770 );
    not g7653 ( n10688 , n22287 );
    nor g7654 ( n22259 , n4168 , n5975 );
    xnor g7655 ( n4228 , n5347 , n31139 );
    xnor g7656 ( n12196 , n21479 , n21842 );
    not g7657 ( n6944 , n19585 );
    xnor g7658 ( n19237 , n932 , n28192 );
    and g7659 ( n2695 , n1604 , n9987 );
    or g7660 ( n12829 , n12474 , n22875 );
    xnor g7661 ( n4620 , n22213 , n25759 );
    and g7662 ( n6308 , n5357 , n1227 );
    not g7663 ( n18370 , n4154 );
    not g7664 ( n25217 , n14441 );
    not g7665 ( n16531 , n27166 );
    not g7666 ( n15181 , n30426 );
    not g7667 ( n7562 , n14434 );
    or g7668 ( n2038 , n23324 , n9178 );
    or g7669 ( n31296 , n26245 , n4327 );
    not g7670 ( n26787 , n3907 );
    not g7671 ( n87 , n14542 );
    and g7672 ( n27837 , n15354 , n31572 );
    and g7673 ( n229 , n13995 , n28550 );
    and g7674 ( n17663 , n5287 , n29228 );
    or g7675 ( n1989 , n872 , n23482 );
    or g7676 ( n1666 , n30178 , n3562 );
    not g7677 ( n5050 , n15993 );
    or g7678 ( n20689 , n7754 , n7792 );
    xnor g7679 ( n21494 , n28175 , n1995 );
    and g7680 ( n13013 , n11844 , n19627 );
    xnor g7681 ( n2288 , n21696 , n29380 );
    or g7682 ( n2077 , n19526 , n25852 );
    and g7683 ( n6228 , n22 , n18471 );
    or g7684 ( n26013 , n12878 , n9419 );
    not g7685 ( n19167 , n16418 );
    xnor g7686 ( n11585 , n24993 , n24391 );
    xnor g7687 ( n17358 , n15510 , n10071 );
    or g7688 ( n28526 , n10867 , n24685 );
    or g7689 ( n22535 , n22756 , n15121 );
    or g7690 ( n11107 , n25488 , n526 );
    not g7691 ( n15884 , n18735 );
    not g7692 ( n18605 , n5306 );
    and g7693 ( n23696 , n14531 , n17528 );
    not g7694 ( n9548 , n25035 );
    not g7695 ( n22916 , n23588 );
    not g7696 ( n28504 , n7651 );
    and g7697 ( n4721 , n2745 , n26617 );
    not g7698 ( n13733 , n534 );
    and g7699 ( n15856 , n30039 , n5219 );
    or g7700 ( n19380 , n25627 , n11305 );
    not g7701 ( n31546 , n24503 );
    xnor g7702 ( n30660 , n3481 , n25276 );
    xnor g7703 ( n4296 , n25527 , n17302 );
    not g7704 ( n16922 , n28452 );
    not g7705 ( n3659 , n30636 );
    nor g7706 ( n12965 , n29923 , n17007 );
    xnor g7707 ( n15753 , n12460 , n31996 );
    not g7708 ( n27367 , n7225 );
    nor g7709 ( n23361 , n14669 , n22814 );
    not g7710 ( n679 , n13145 );
    and g7711 ( n28902 , n30463 , n16172 );
    or g7712 ( n18297 , n2207 , n15459 );
    and g7713 ( n12820 , n12474 , n2112 );
    or g7714 ( n26582 , n15251 , n12254 );
    xnor g7715 ( n10925 , n20312 , n31394 );
    nor g7716 ( n9740 , n6940 , n26200 );
    xnor g7717 ( n23142 , n25988 , n6755 );
    or g7718 ( n24718 , n5492 , n3098 );
    xnor g7719 ( n31998 , n8999 , n25527 );
    xnor g7720 ( n24448 , n23659 , n21268 );
    and g7721 ( n23192 , n4932 , n25961 );
    and g7722 ( n5615 , n24240 , n9465 );
    not g7723 ( n28809 , n31702 );
    or g7724 ( n10424 , n30769 , n29665 );
    xnor g7725 ( n9205 , n10759 , n31168 );
    xnor g7726 ( n27477 , n24637 , n8267 );
    not g7727 ( n20959 , n921 );
    not g7728 ( n8317 , n2589 );
    or g7729 ( n30261 , n27522 , n376 );
    not g7730 ( n20093 , n13482 );
    not g7731 ( n23226 , n530 );
    xnor g7732 ( n2071 , n14031 , n18167 );
    nor g7733 ( n23859 , n11711 , n31856 );
    xnor g7734 ( n19805 , n20190 , n20404 );
    buf g7735 ( n8987 , n16384 );
    and g7736 ( n31243 , n12985 , n9218 );
    not g7737 ( n16168 , n26300 );
    nor g7738 ( n267 , n19538 , n13859 );
    not g7739 ( n19291 , n2533 );
    not g7740 ( n14274 , n22850 );
    not g7741 ( n30771 , n9310 );
    xnor g7742 ( n15006 , n26017 , n19743 );
    or g7743 ( n24736 , n16702 , n4136 );
    xnor g7744 ( n21017 , n10837 , n11361 );
    xnor g7745 ( n10912 , n30514 , n24066 );
    xor g7746 ( n29478 , n10272 , n8161 );
    not g7747 ( n17840 , n5332 );
    or g7748 ( n20406 , n26820 , n31560 );
    not g7749 ( n16946 , n8654 );
    or g7750 ( n15657 , n9540 , n6422 );
    and g7751 ( n15025 , n19184 , n13703 );
    nor g7752 ( n9181 , n13264 , n22577 );
    or g7753 ( n15882 , n12556 , n1691 );
    not g7754 ( n28778 , n23772 );
    or g7755 ( n30573 , n21357 , n7410 );
    or g7756 ( n1735 , n29571 , n13464 );
    xnor g7757 ( n13234 , n12822 , n13963 );
    xnor g7758 ( n5915 , n20402 , n11555 );
    xnor g7759 ( n22819 , n27903 , n27414 );
    not g7760 ( n8924 , n31032 );
    not g7761 ( n3656 , n14036 );
    and g7762 ( n26923 , n11514 , n671 );
    and g7763 ( n22209 , n26413 , n9591 );
    not g7764 ( n2302 , n26192 );
    not g7765 ( n24681 , n1307 );
    xnor g7766 ( n2177 , n7389 , n1813 );
    not g7767 ( n11698 , n28983 );
    and g7768 ( n13747 , n5117 , n28344 );
    or g7769 ( n10418 , n17934 , n16761 );
    xnor g7770 ( n7905 , n23088 , n6957 );
    xnor g7771 ( n1700 , n30596 , n19525 );
    nor g7772 ( n28070 , n26337 , n14649 );
    xnor g7773 ( n5793 , n1950 , n5443 );
    or g7774 ( n3356 , n22244 , n20848 );
    not g7775 ( n2877 , n6493 );
    xnor g7776 ( n18209 , n2925 , n25805 );
    not g7777 ( n26265 , n22184 );
    xnor g7778 ( n12139 , n30563 , n8688 );
    not g7779 ( n12190 , n1670 );
    xnor g7780 ( n476 , n29141 , n11035 );
    not g7781 ( n18474 , n25320 );
    or g7782 ( n21031 , n8111 , n10315 );
    not g7783 ( n20964 , n29659 );
    xnor g7784 ( n804 , n16130 , n16701 );
    not g7785 ( n31486 , n25786 );
    and g7786 ( n10873 , n10604 , n644 );
    and g7787 ( n16849 , n30778 , n17994 );
    xnor g7788 ( n22029 , n26410 , n10524 );
    xnor g7789 ( n17596 , n10256 , n15400 );
    not g7790 ( n3197 , n29661 );
    not g7791 ( n1199 , n21712 );
    not g7792 ( n27723 , n2150 );
    nor g7793 ( n6831 , n29052 , n16092 );
    xnor g7794 ( n2147 , n9546 , n15077 );
    not g7795 ( n487 , n29346 );
    not g7796 ( n11987 , n25493 );
    and g7797 ( n3615 , n31912 , n28557 );
    xor g7798 ( n24775 , n31116 , n28734 );
    or g7799 ( n12591 , n18779 , n29260 );
    and g7800 ( n164 , n18091 , n23331 );
    or g7801 ( n3204 , n32000 , n1101 );
    or g7802 ( n13956 , n28720 , n16599 );
    nor g7803 ( n15824 , n22345 , n19358 );
    not g7804 ( n22697 , n28772 );
    or g7805 ( n5918 , n23846 , n22271 );
    or g7806 ( n14022 , n14750 , n24663 );
    or g7807 ( n27915 , n15129 , n24427 );
    nor g7808 ( n30129 , n2568 , n14708 );
    nor g7809 ( n22944 , n18518 , n17645 );
    xnor g7810 ( n13385 , n10294 , n23530 );
    not g7811 ( n9931 , n8638 );
    and g7812 ( n9556 , n2541 , n31365 );
    buf g7813 ( n22139 , n10255 );
    not g7814 ( n3875 , n16835 );
    or g7815 ( n31047 , n17257 , n3829 );
    or g7816 ( n27053 , n15495 , n30901 );
    or g7817 ( n23036 , n20276 , n28173 );
    and g7818 ( n30849 , n6443 , n2084 );
    and g7819 ( n14218 , n12529 , n17181 );
    and g7820 ( n9798 , n7446 , n25319 );
    not g7821 ( n20267 , n3810 );
    nor g7822 ( n26662 , n26156 , n10168 );
    xnor g7823 ( n11735 , n11704 , n20967 );
    and g7824 ( n32019 , n31461 , n13756 );
    and g7825 ( n1504 , n9042 , n13911 );
    not g7826 ( n15361 , n12827 );
    and g7827 ( n2233 , n28941 , n29953 );
    and g7828 ( n25528 , n9597 , n10457 );
    or g7829 ( n24312 , n19756 , n5100 );
    xnor g7830 ( n22315 , n18941 , n8023 );
    or g7831 ( n17806 , n30270 , n17339 );
    and g7832 ( n7136 , n30737 , n24103 );
    xnor g7833 ( n17103 , n23133 , n17585 );
    not g7834 ( n25675 , n9537 );
    or g7835 ( n31275 , n7970 , n9298 );
    nor g7836 ( n2187 , n15588 , n24837 );
    nor g7837 ( n29011 , n20273 , n15529 );
    not g7838 ( n5480 , n26072 );
    or g7839 ( n14322 , n29262 , n13771 );
    and g7840 ( n29081 , n11633 , n9450 );
    and g7841 ( n16550 , n18081 , n6019 );
    xnor g7842 ( n5382 , n28927 , n6717 );
    nor g7843 ( n29040 , n23842 , n12739 );
    or g7844 ( n10022 , n29005 , n25795 );
    or g7845 ( n4301 , n28223 , n15386 );
    xnor g7846 ( n20212 , n25990 , n12554 );
    xor g7847 ( n3352 , n16518 , n23182 );
    xnor g7848 ( n30951 , n6884 , n25211 );
    or g7849 ( n19402 , n2915 , n17610 );
    not g7850 ( n14388 , n1748 );
    xnor g7851 ( n31830 , n16710 , n17615 );
    and g7852 ( n3308 , n14971 , n29815 );
    and g7853 ( n9129 , n19952 , n20201 );
    xnor g7854 ( n30900 , n30751 , n24219 );
    or g7855 ( n727 , n16592 , n10480 );
    not g7856 ( n20604 , n27045 );
    not g7857 ( n27117 , n7778 );
    xnor g7858 ( n29309 , n3319 , n18743 );
    xnor g7859 ( n31785 , n12267 , n650 );
    not g7860 ( n27334 , n3449 );
    xnor g7861 ( n7304 , n25044 , n30540 );
    and g7862 ( n24417 , n29501 , n23478 );
    or g7863 ( n30008 , n10094 , n6642 );
    not g7864 ( n15837 , n1952 );
    nor g7865 ( n16921 , n17305 , n10538 );
    xnor g7866 ( n23685 , n30167 , n31301 );
    nor g7867 ( n7261 , n23079 , n11908 );
    xnor g7868 ( n21723 , n2651 , n17358 );
    nor g7869 ( n156 , n2702 , n17623 );
    xnor g7870 ( n4077 , n1209 , n2848 );
    not g7871 ( n6900 , n16420 );
    and g7872 ( n11910 , n15931 , n7114 );
    xnor g7873 ( n1318 , n19977 , n12776 );
    nor g7874 ( n21270 , n13075 , n13348 );
    and g7875 ( n12100 , n24279 , n19265 );
    or g7876 ( n14279 , n19695 , n6386 );
    not g7877 ( n13548 , n18370 );
    and g7878 ( n22636 , n31550 , n27871 );
    xnor g7879 ( n8305 , n6757 , n27859 );
    xnor g7880 ( n6655 , n25061 , n20449 );
    nor g7881 ( n25516 , n1570 , n20642 );
    nor g7882 ( n21205 , n22244 , n31049 );
    xnor g7883 ( n9705 , n2939 , n2231 );
    xnor g7884 ( n18374 , n29131 , n4433 );
    xnor g7885 ( n13961 , n9237 , n20602 );
    or g7886 ( n25202 , n31053 , n4873 );
    xnor g7887 ( n28938 , n16075 , n14106 );
    not g7888 ( n6896 , n12998 );
    not g7889 ( n10717 , n23523 );
    not g7890 ( n555 , n17615 );
    nor g7891 ( n9326 , n26959 , n23511 );
    not g7892 ( n30896 , n24596 );
    not g7893 ( n24741 , n22433 );
    xnor g7894 ( n1776 , n22468 , n3591 );
    and g7895 ( n30154 , n16696 , n30076 );
    xnor g7896 ( n29710 , n24809 , n24682 );
    not g7897 ( n4264 , n22845 );
    nor g7898 ( n29771 , n31481 , n13859 );
    or g7899 ( n26597 , n27805 , n27008 );
    and g7900 ( n2273 , n31255 , n19133 );
    not g7901 ( n22938 , n18725 );
    not g7902 ( n31884 , n11177 );
    xnor g7903 ( n21265 , n29311 , n1898 );
    and g7904 ( n4467 , n8749 , n19416 );
    xor g7905 ( n21773 , n12397 , n29515 );
    or g7906 ( n3424 , n22045 , n2943 );
    or g7907 ( n15378 , n5527 , n27293 );
    not g7908 ( n14481 , n16972 );
    not g7909 ( n3067 , n12128 );
    xnor g7910 ( n12271 , n15106 , n14718 );
    not g7911 ( n7013 , n30096 );
    not g7912 ( n13795 , n16967 );
    nor g7913 ( n18771 , n255 , n21777 );
    not g7914 ( n25838 , n9842 );
    and g7915 ( n18999 , n15194 , n25123 );
    xnor g7916 ( n25429 , n27885 , n12920 );
    or g7917 ( n17340 , n2887 , n8541 );
    and g7918 ( n30712 , n15285 , n20685 );
    not g7919 ( n7495 , n5622 );
    or g7920 ( n19794 , n13514 , n31193 );
    not g7921 ( n22413 , n31362 );
    or g7922 ( n11448 , n28986 , n21586 );
    nor g7923 ( n18553 , n30067 , n9338 );
    nor g7924 ( n21146 , n4213 , n31604 );
    and g7925 ( n28275 , n31219 , n4265 );
    and g7926 ( n13093 , n30835 , n23793 );
    or g7927 ( n10402 , n18967 , n22484 );
    or g7928 ( n21199 , n3788 , n16263 );
    or g7929 ( n10678 , n3166 , n28869 );
    and g7930 ( n10591 , n17400 , n17989 );
    nor g7931 ( n6233 , n4332 , n25398 );
    and g7932 ( n23492 , n7544 , n27096 );
    xnor g7933 ( n16858 , n28469 , n27380 );
    and g7934 ( n3961 , n12834 , n17408 );
    nor g7935 ( n10021 , n23829 , n13363 );
    not g7936 ( n8815 , n23639 );
    xnor g7937 ( n8404 , n7209 , n31722 );
    and g7938 ( n750 , n4290 , n918 );
    or g7939 ( n5657 , n13252 , n19831 );
    or g7940 ( n7003 , n9682 , n6731 );
    xnor g7941 ( n17677 , n22917 , n23960 );
    not g7942 ( n461 , n25596 );
    xnor g7943 ( n18936 , n14465 , n28389 );
    and g7944 ( n1595 , n5601 , n5495 );
    not g7945 ( n18193 , n23914 );
    buf g7946 ( n13549 , n19080 );
    not g7947 ( n29817 , n20192 );
    and g7948 ( n2149 , n19632 , n18667 );
    xnor g7949 ( n17990 , n30839 , n6646 );
    xnor g7950 ( n20844 , n24644 , n13563 );
    not g7951 ( n23675 , n6188 );
    or g7952 ( n10235 , n3765 , n10315 );
    or g7953 ( n7286 , n21525 , n8133 );
    not g7954 ( n25882 , n30061 );
    not g7955 ( n19834 , n4248 );
    not g7956 ( n11301 , n12601 );
    or g7957 ( n22589 , n23848 , n4606 );
    xnor g7958 ( n29720 , n7829 , n5112 );
    and g7959 ( n28276 , n27588 , n13368 );
    not g7960 ( n22429 , n25373 );
    not g7961 ( n30504 , n8356 );
    xor g7962 ( n11425 , n5172 , n14992 );
    not g7963 ( n26720 , n5541 );
    and g7964 ( n13866 , n26219 , n16105 );
    or g7965 ( n9230 , n22905 , n20687 );
    not g7966 ( n27155 , n29248 );
    not g7967 ( n26176 , n26695 );
    not g7968 ( n7709 , n30165 );
    xnor g7969 ( n15782 , n16209 , n28638 );
    not g7970 ( n23022 , n24643 );
    xnor g7971 ( n10846 , n12145 , n16113 );
    not g7972 ( n1317 , n27 );
    xnor g7973 ( n1210 , n351 , n25515 );
    not g7974 ( n11626 , n15878 );
    nor g7975 ( n22274 , n8714 , n22489 );
    and g7976 ( n1187 , n11395 , n9212 );
    not g7977 ( n9463 , n1667 );
    and g7978 ( n29900 , n21040 , n28994 );
    xnor g7979 ( n24536 , n29097 , n11459 );
    or g7980 ( n12662 , n24429 , n20871 );
    xnor g7981 ( n4194 , n174 , n20501 );
    nor g7982 ( n4575 , n13204 , n5731 );
    not g7983 ( n4999 , n8624 );
    xnor g7984 ( n26747 , n25119 , n14205 );
    not g7985 ( n8921 , n16152 );
    and g7986 ( n12701 , n9046 , n1373 );
    xnor g7987 ( n9717 , n5407 , n31101 );
    or g7988 ( n19073 , n21912 , n24337 );
    or g7989 ( n11772 , n29156 , n22188 );
    not g7990 ( n31497 , n7604 );
    xnor g7991 ( n30273 , n25619 , n17082 );
    or g7992 ( n24821 , n6713 , n5780 );
    and g7993 ( n10224 , n31065 , n3549 );
    and g7994 ( n5369 , n24632 , n23273 );
    xnor g7995 ( n22623 , n2956 , n25616 );
    and g7996 ( n10496 , n15663 , n3591 );
    not g7997 ( n2115 , n19572 );
    or g7998 ( n3583 , n15987 , n11624 );
    and g7999 ( n8412 , n7393 , n14041 );
    not g8000 ( n4586 , n31295 );
    and g8001 ( n11597 , n8141 , n28403 );
    nor g8002 ( n21175 , n23290 , n7684 );
    or g8003 ( n18073 , n17321 , n309 );
    not g8004 ( n20043 , n30326 );
    xnor g8005 ( n8688 , n8064 , n27848 );
    xnor g8006 ( n5454 , n28983 , n15999 );
    not g8007 ( n29150 , n26969 );
    nor g8008 ( n12345 , n2218 , n11820 );
    and g8009 ( n3329 , n1506 , n17921 );
    or g8010 ( n29002 , n4534 , n30583 );
    and g8011 ( n4146 , n29130 , n19104 );
    not g8012 ( n25626 , n26362 );
    not g8013 ( n20906 , n10981 );
    xnor g8014 ( n30083 , n24130 , n23646 );
    or g8015 ( n25780 , n9001 , n3327 );
    xnor g8016 ( n23262 , n20005 , n18072 );
    not g8017 ( n22516 , n20998 );
    xnor g8018 ( n2258 , n6626 , n27805 );
    or g8019 ( n15508 , n26894 , n19693 );
    not g8020 ( n25510 , n3869 );
    not g8021 ( n25862 , n5453 );
    not g8022 ( n21535 , n11745 );
    xnor g8023 ( n753 , n18972 , n3307 );
    nor g8024 ( n25571 , n24988 , n14798 );
    not g8025 ( n21308 , n28638 );
    not g8026 ( n11858 , n12169 );
    xnor g8027 ( n17879 , n23306 , n9653 );
    not g8028 ( n5281 , n1635 );
    and g8029 ( n17280 , n20458 , n16018 );
    and g8030 ( n9423 , n2591 , n14867 );
    xnor g8031 ( n550 , n19297 , n17293 );
    or g8032 ( n22588 , n22558 , n873 );
    and g8033 ( n12268 , n6194 , n8907 );
    not g8034 ( n16418 , n894 );
    and g8035 ( n5463 , n2114 , n17202 );
    nor g8036 ( n6151 , n10400 , n30089 );
    not g8037 ( n6757 , n17900 );
    not g8038 ( n21995 , n28006 );
    xnor g8039 ( n26226 , n15334 , n8584 );
    and g8040 ( n31749 , n23969 , n8741 );
    nor g8041 ( n21094 , n12140 , n17289 );
    and g8042 ( n20451 , n26753 , n20583 );
    not g8043 ( n29782 , n14186 );
    or g8044 ( n11758 , n3490 , n2811 );
    nor g8045 ( n30848 , n16778 , n1688 );
    or g8046 ( n11518 , n11348 , n2076 );
    xnor g8047 ( n9578 , n13613 , n16801 );
    xnor g8048 ( n17159 , n8667 , n3401 );
    xnor g8049 ( n23714 , n28654 , n27531 );
    not g8050 ( n12111 , n30176 );
    nor g8051 ( n3681 , n12138 , n16559 );
    and g8052 ( n24764 , n17029 , n29656 );
    or g8053 ( n22419 , n12992 , n11478 );
    and g8054 ( n27437 , n3074 , n199 );
    nor g8055 ( n15916 , n4175 , n10847 );
    xnor g8056 ( n10842 , n7348 , n3076 );
    or g8057 ( n31978 , n16279 , n28716 );
    not g8058 ( n2339 , n21643 );
    or g8059 ( n18571 , n7658 , n19743 );
    or g8060 ( n28321 , n6295 , n5098 );
    or g8061 ( n11536 , n20365 , n18595 );
    xnor g8062 ( n8627 , n10155 , n28034 );
    not g8063 ( n29143 , n18448 );
    not g8064 ( n23871 , n4561 );
    and g8065 ( n25615 , n2952 , n13590 );
    or g8066 ( n26770 , n13975 , n29770 );
    not g8067 ( n568 , n18997 );
    not g8068 ( n27459 , n4120 );
    nor g8069 ( n23314 , n14872 , n19643 );
    and g8070 ( n30752 , n22051 , n31731 );
    not g8071 ( n1484 , n14464 );
    xor g8072 ( n8669 , n14755 , n16110 );
    and g8073 ( n8277 , n22873 , n9355 );
    xnor g8074 ( n23901 , n3858 , n6626 );
    xnor g8075 ( n10077 , n2425 , n27023 );
    and g8076 ( n1990 , n18986 , n7444 );
    or g8077 ( n5357 , n10739 , n7018 );
    not g8078 ( n434 , n13677 );
    xnor g8079 ( n7657 , n25821 , n5496 );
    nor g8080 ( n32002 , n24184 , n29059 );
    xnor g8081 ( n23649 , n24183 , n16163 );
    and g8082 ( n23743 , n11358 , n29273 );
    and g8083 ( n31788 , n25445 , n29668 );
    not g8084 ( n23518 , n17843 );
    not g8085 ( n14443 , n31231 );
    xnor g8086 ( n12004 , n3351 , n26319 );
    not g8087 ( n12958 , n16054 );
    or g8088 ( n1836 , n3758 , n21785 );
    or g8089 ( n19543 , n387 , n20227 );
    or g8090 ( n15766 , n30600 , n10025 );
    not g8091 ( n7582 , n29119 );
    xnor g8092 ( n26844 , n1342 , n29901 );
    xnor g8093 ( n18278 , n21305 , n9034 );
    or g8094 ( n21207 , n21755 , n10572 );
    or g8095 ( n21923 , n29000 , n22614 );
    not g8096 ( n14700 , n25272 );
    not g8097 ( n22573 , n24471 );
    buf g8098 ( n26117 , n31757 );
    xnor g8099 ( n169 , n14121 , n21603 );
    not g8100 ( n17537 , n12232 );
    not g8101 ( n15210 , n11387 );
    and g8102 ( n14919 , n3380 , n3026 );
    or g8103 ( n17064 , n4213 , n28103 );
    xnor g8104 ( n24202 , n21328 , n13263 );
    or g8105 ( n22354 , n1887 , n29272 );
    or g8106 ( n15903 , n16620 , n30093 );
    xnor g8107 ( n4727 , n23743 , n730 );
    and g8108 ( n26129 , n30353 , n14060 );
    xnor g8109 ( n6641 , n24054 , n27177 );
    xnor g8110 ( n13785 , n31926 , n30904 );
    or g8111 ( n3958 , n12064 , n8073 );
    not g8112 ( n28256 , n17205 );
    not g8113 ( n9328 , n15100 );
    and g8114 ( n24956 , n14286 , n24988 );
    not g8115 ( n6130 , n15981 );
    and g8116 ( n11854 , n9007 , n7286 );
    xnor g8117 ( n2714 , n29635 , n4539 );
    not g8118 ( n12513 , n20251 );
    or g8119 ( n13001 , n7201 , n26539 );
    or g8120 ( n10211 , n23469 , n4862 );
    or g8121 ( n24079 , n18452 , n22184 );
    or g8122 ( n31148 , n4817 , n22335 );
    not g8123 ( n20690 , n14123 );
    xnor g8124 ( n31614 , n3036 , n31204 );
    xnor g8125 ( n30968 , n14690 , n3307 );
    and g8126 ( n29178 , n31607 , n19461 );
    and g8127 ( n11058 , n26208 , n24 );
    not g8128 ( n13313 , n10730 );
    not g8129 ( n6287 , n18850 );
    and g8130 ( n28880 , n27344 , n22974 );
    or g8131 ( n21675 , n27374 , n9638 );
    nor g8132 ( n1017 , n24630 , n10841 );
    xnor g8133 ( n26298 , n1237 , n21237 );
    and g8134 ( n18468 , n4718 , n29573 );
    not g8135 ( n9868 , n20541 );
    not g8136 ( n16391 , n27390 );
    or g8137 ( n16332 , n9939 , n6426 );
    nor g8138 ( n473 , n23726 , n23470 );
    not g8139 ( n1275 , n11600 );
    and g8140 ( n18976 , n21494 , n31783 );
    xnor g8141 ( n30489 , n2416 , n24327 );
    not g8142 ( n6674 , n28417 );
    and g8143 ( n14747 , n22907 , n21104 );
    xnor g8144 ( n5739 , n21814 , n30936 );
    xnor g8145 ( n3333 , n7454 , n13933 );
    not g8146 ( n23848 , n18507 );
    not g8147 ( n4414 , n18322 );
    or g8148 ( n19829 , n11734 , n8167 );
    nor g8149 ( n4170 , n17704 , n12880 );
    not g8150 ( n25186 , n26862 );
    not g8151 ( n10152 , n20468 );
    not g8152 ( n5646 , n20279 );
    or g8153 ( n24186 , n12210 , n14936 );
    not g8154 ( n13194 , n9778 );
    nor g8155 ( n3 , n24807 , n20854 );
    not g8156 ( n13766 , n4322 );
    or g8157 ( n7040 , n20304 , n12460 );
    nor g8158 ( n27408 , n27354 , n20334 );
    and g8159 ( n11582 , n17225 , n16217 );
    not g8160 ( n28319 , n25117 );
    nor g8161 ( n16526 , n30887 , n11771 );
    nor g8162 ( n20372 , n1128 , n314 );
    xnor g8163 ( n22766 , n15030 , n30308 );
    and g8164 ( n4323 , n26166 , n7964 );
    and g8165 ( n13531 , n3204 , n24723 );
    nor g8166 ( n26801 , n2483 , n7663 );
    nor g8167 ( n11317 , n15465 , n5726 );
    or g8168 ( n21380 , n16114 , n6328 );
    nor g8169 ( n30604 , n9340 , n2831 );
    or g8170 ( n22014 , n12627 , n28302 );
    and g8171 ( n16429 , n8066 , n26600 );
    or g8172 ( n19868 , n17109 , n15948 );
    not g8173 ( n26959 , n2802 );
    or g8174 ( n6461 , n10832 , n27735 );
    or g8175 ( n19175 , n27108 , n24411 );
    not g8176 ( n21253 , n2678 );
    xnor g8177 ( n31563 , n5257 , n10574 );
    not g8178 ( n16189 , n9635 );
    xnor g8179 ( n29939 , n763 , n4393 );
    or g8180 ( n27894 , n20729 , n26628 );
    or g8181 ( n12589 , n5109 , n9994 );
    nor g8182 ( n3457 , n7665 , n10770 );
    not g8183 ( n8819 , n20131 );
    not g8184 ( n6539 , n22707 );
    or g8185 ( n17989 , n4608 , n30552 );
    xor g8186 ( n31679 , n30274 , n15191 );
    or g8187 ( n29621 , n1721 , n16955 );
    and g8188 ( n16854 , n1460 , n26682 );
    xor g8189 ( n3461 , n4045 , n21200 );
    not g8190 ( n14640 , n8394 );
    xnor g8191 ( n23968 , n7627 , n2840 );
    or g8192 ( n12847 , n2852 , n4242 );
    and g8193 ( n27290 , n14459 , n8740 );
    and g8194 ( n11038 , n3503 , n65 );
    buf g8195 ( n27538 , n21921 );
    or g8196 ( n27417 , n14899 , n30518 );
    and g8197 ( n31715 , n12006 , n7418 );
    or g8198 ( n3652 , n7024 , n27484 );
    not g8199 ( n23468 , n23533 );
    not g8200 ( n12284 , n2885 );
    not g8201 ( n1205 , n22280 );
    xnor g8202 ( n27565 , n2918 , n26665 );
    xnor g8203 ( n7313 , n26714 , n23104 );
    or g8204 ( n30911 , n17089 , n4393 );
    nor g8205 ( n14811 , n24418 , n31843 );
    and g8206 ( n17512 , n12107 , n30762 );
    not g8207 ( n22020 , n23928 );
    and g8208 ( n21430 , n25697 , n22668 );
    xnor g8209 ( n31869 , n13054 , n27901 );
    or g8210 ( n15881 , n23705 , n14122 );
    xnor g8211 ( n22016 , n9242 , n23254 );
    not g8212 ( n15118 , n18113 );
    xnor g8213 ( n8685 , n7602 , n1434 );
    not g8214 ( n10452 , n14423 );
    and g8215 ( n20955 , n16576 , n19580 );
    xnor g8216 ( n16365 , n17343 , n13950 );
    nor g8217 ( n4197 , n30607 , n19050 );
    not g8218 ( n11507 , n876 );
    or g8219 ( n18962 , n24196 , n20958 );
    xnor g8220 ( n16264 , n24760 , n5315 );
    buf g8221 ( n21050 , n25306 );
    not g8222 ( n29920 , n10350 );
    xnor g8223 ( n12116 , n2595 , n15436 );
    xnor g8224 ( n27625 , n18385 , n31725 );
    not g8225 ( n20055 , n15517 );
    xnor g8226 ( n16487 , n13650 , n12017 );
    xnor g8227 ( n18381 , n10652 , n632 );
    xnor g8228 ( n21343 , n11214 , n532 );
    not g8229 ( n30758 , n11008 );
    and g8230 ( n23234 , n30764 , n5093 );
    xor g8231 ( n21890 , n6414 , n20066 );
    not g8232 ( n2263 , n28843 );
    xnor g8233 ( n10615 , n22883 , n26595 );
    xor g8234 ( n6789 , n27520 , n18667 );
    xnor g8235 ( n13016 , n8580 , n10713 );
    xnor g8236 ( n14277 , n19862 , n2290 );
    xnor g8237 ( n25204 , n2923 , n16260 );
    xnor g8238 ( n4190 , n16063 , n583 );
    xnor g8239 ( n25300 , n19672 , n9661 );
    not g8240 ( n27992 , n442 );
    xnor g8241 ( n19621 , n8057 , n10599 );
    xnor g8242 ( n14988 , n7548 , n2665 );
    nor g8243 ( n26716 , n2722 , n30414 );
    and g8244 ( n18533 , n21537 , n10014 );
    not g8245 ( n29641 , n1066 );
    not g8246 ( n1665 , n3911 );
    not g8247 ( n8597 , n13726 );
    xnor g8248 ( n16163 , n8561 , n31727 );
    xnor g8249 ( n12562 , n26867 , n14828 );
    not g8250 ( n1450 , n5792 );
    or g8251 ( n10953 , n30227 , n6384 );
    or g8252 ( n30222 , n30943 , n23735 );
    and g8253 ( n27628 , n27999 , n12000 );
    or g8254 ( n28917 , n14831 , n7940 );
    or g8255 ( n19430 , n15118 , n6798 );
    xnor g8256 ( n4403 , n20924 , n4048 );
    nor g8257 ( n12654 , n8150 , n7644 );
    and g8258 ( n14815 , n6532 , n23780 );
    or g8259 ( n16618 , n26929 , n4926 );
    xnor g8260 ( n29740 , n27885 , n11065 );
    and g8261 ( n12588 , n20484 , n7776 );
    xnor g8262 ( n17180 , n10571 , n6383 );
    nor g8263 ( n25859 , n17019 , n9263 );
    or g8264 ( n15908 , n16799 , n27135 );
    not g8265 ( n1322 , n10350 );
    not g8266 ( n594 , n19066 );
    and g8267 ( n7505 , n1081 , n30773 );
    not g8268 ( n31257 , n13148 );
    xnor g8269 ( n29836 , n8527 , n15846 );
    and g8270 ( n25461 , n6836 , n5559 );
    xnor g8271 ( n18170 , n10345 , n12204 );
    xnor g8272 ( n27882 , n11827 , n10325 );
    nor g8273 ( n1049 , n6125 , n15716 );
    xnor g8274 ( n8806 , n6758 , n13116 );
    not g8275 ( n10287 , n14106 );
    or g8276 ( n8227 , n23676 , n16508 );
    not g8277 ( n3011 , n20836 );
    not g8278 ( n29688 , n24977 );
    or g8279 ( n10160 , n31184 , n24606 );
    or g8280 ( n12452 , n25457 , n23864 );
    xor g8281 ( n28632 , n24704 , n6488 );
    xnor g8282 ( n13315 , n29544 , n11346 );
    xor g8283 ( n17298 , n21437 , n4315 );
    not g8284 ( n3464 , n3849 );
    or g8285 ( n3825 , n24715 , n20855 );
    and g8286 ( n29204 , n23821 , n703 );
    nor g8287 ( n3216 , n13137 , n18990 );
    xnor g8288 ( n19987 , n21668 , n23453 );
    or g8289 ( n23733 , n29709 , n12525 );
    not g8290 ( n14248 , n7011 );
    or g8291 ( n11084 , n17542 , n31294 );
    and g8292 ( n22693 , n18704 , n10099 );
    or g8293 ( n28888 , n28397 , n9321 );
    xnor g8294 ( n28289 , n28980 , n31453 );
    or g8295 ( n26554 , n30561 , n4283 );
    xnor g8296 ( n3534 , n28057 , n17867 );
    not g8297 ( n25299 , n6636 );
    or g8298 ( n15659 , n4158 , n17210 );
    nor g8299 ( n463 , n15502 , n30030 );
    nor g8300 ( n9791 , n2660 , n13247 );
    nor g8301 ( n12795 , n3614 , n20583 );
    nor g8302 ( n17035 , n1250 , n2724 );
    or g8303 ( n19314 , n21603 , n17819 );
    and g8304 ( n4640 , n28222 , n22451 );
    and g8305 ( n6398 , n29180 , n5869 );
    and g8306 ( n17488 , n4910 , n1942 );
    nor g8307 ( n26084 , n632 , n3655 );
    not g8308 ( n21160 , n20153 );
    xnor g8309 ( n7192 , n8347 , n27083 );
    or g8310 ( n29628 , n2888 , n20044 );
    and g8311 ( n30015 , n410 , n22932 );
    nor g8312 ( n24229 , n21466 , n22157 );
    or g8313 ( n17403 , n28324 , n31775 );
    or g8314 ( n8810 , n7697 , n24203 );
    not g8315 ( n4507 , n9684 );
    xnor g8316 ( n172 , n28158 , n22393 );
    not g8317 ( n1724 , n3676 );
    not g8318 ( n20536 , n10158 );
    not g8319 ( n7636 , n26560 );
    or g8320 ( n5445 , n9124 , n19186 );
    not g8321 ( n1004 , n14136 );
    not g8322 ( n8278 , n13572 );
    not g8323 ( n12074 , n6867 );
    and g8324 ( n11285 , n23267 , n21051 );
    not g8325 ( n13011 , n2232 );
    or g8326 ( n6341 , n23071 , n1444 );
    or g8327 ( n11055 , n9220 , n29654 );
    or g8328 ( n7428 , n10721 , n1102 );
    xnor g8329 ( n4169 , n16674 , n11610 );
    nor g8330 ( n31469 , n13262 , n12794 );
    nor g8331 ( n10308 , n15358 , n17832 );
    not g8332 ( n7902 , n19090 );
    or g8333 ( n11930 , n31782 , n22301 );
    xnor g8334 ( n18870 , n9468 , n11072 );
    not g8335 ( n5719 , n9888 );
    xnor g8336 ( n8108 , n18450 , n10737 );
    not g8337 ( n205 , n19654 );
    not g8338 ( n5352 , n31491 );
    nor g8339 ( n21755 , n5895 , n2749 );
    and g8340 ( n29927 , n6155 , n12010 );
    xnor g8341 ( n21349 , n4299 , n17798 );
    nor g8342 ( n29603 , n1873 , n10382 );
    or g8343 ( n24162 , n20453 , n8763 );
    not g8344 ( n3377 , n6381 );
    and g8345 ( n12267 , n19063 , n3045 );
    xnor g8346 ( n2072 , n24933 , n25453 );
    xnor g8347 ( n8770 , n16730 , n25826 );
    not g8348 ( n22915 , n10943 );
    nor g8349 ( n8171 , n26328 , n8612 );
    or g8350 ( n12930 , n30305 , n4529 );
    xnor g8351 ( n28593 , n314 , n26385 );
    not g8352 ( n16266 , n7676 );
    xnor g8353 ( n10633 , n7244 , n6349 );
    not g8354 ( n29793 , n5816 );
    or g8355 ( n20950 , n13236 , n19657 );
    xnor g8356 ( n30228 , n3998 , n10687 );
    xor g8357 ( n9193 , n9365 , n1416 );
    not g8358 ( n26078 , n20116 );
    nor g8359 ( n21256 , n13210 , n25913 );
    and g8360 ( n28448 , n12498 , n19055 );
    xnor g8361 ( n21850 , n22657 , n7593 );
    not g8362 ( n26032 , n16200 );
    xnor g8363 ( n14445 , n25704 , n21960 );
    xnor g8364 ( n23407 , n6433 , n29533 );
    xor g8365 ( n2360 , n18710 , n1669 );
    not g8366 ( n8827 , n19405 );
    nor g8367 ( n11315 , n7354 , n4277 );
    xnor g8368 ( n25366 , n26935 , n9883 );
    not g8369 ( n15066 , n14361 );
    or g8370 ( n2031 , n4930 , n6748 );
    not g8371 ( n20388 , n10619 );
    not g8372 ( n12460 , n1102 );
    and g8373 ( n22220 , n21309 , n30571 );
    not g8374 ( n14924 , n24405 );
    or g8375 ( n29537 , n21205 , n14053 );
    xnor g8376 ( n21209 , n20597 , n3711 );
    and g8377 ( n12626 , n15347 , n13153 );
    not g8378 ( n2251 , n28281 );
    or g8379 ( n24616 , n25991 , n679 );
    not g8380 ( n23101 , n30419 );
    or g8381 ( n26538 , n20565 , n9219 );
    or g8382 ( n30773 , n29851 , n12827 );
    nor g8383 ( n9838 , n21492 , n14646 );
    not g8384 ( n3649 , n18148 );
    or g8385 ( n25744 , n19985 , n5285 );
    xnor g8386 ( n17751 , n25946 , n29654 );
    not g8387 ( n17270 , n8732 );
    not g8388 ( n31239 , n11834 );
    or g8389 ( n18340 , n31006 , n18285 );
    not g8390 ( n11015 , n20448 );
    and g8391 ( n31084 , n16159 , n11409 );
    xnor g8392 ( n9746 , n31807 , n5018 );
    not g8393 ( n23660 , n12251 );
    not g8394 ( n21731 , n1979 );
    xnor g8395 ( n8841 , n757 , n20881 );
    and g8396 ( n23691 , n22883 , n20001 );
    nor g8397 ( n28820 , n26607 , n7946 );
    xnor g8398 ( n18382 , n12625 , n14954 );
    xnor g8399 ( n15476 , n23285 , n14013 );
    or g8400 ( n31911 , n12054 , n22774 );
    or g8401 ( n4064 , n24016 , n16014 );
    not g8402 ( n9840 , n9163 );
    xnor g8403 ( n2910 , n1651 , n21504 );
    not g8404 ( n12978 , n12055 );
    xnor g8405 ( n575 , n6002 , n31725 );
    xnor g8406 ( n30622 , n1714 , n31735 );
    or g8407 ( n11657 , n22895 , n5450 );
    not g8408 ( n16675 , n16202 );
    not g8409 ( n22226 , n28627 );
    not g8410 ( n24600 , n28256 );
    or g8411 ( n20102 , n944 , n23546 );
    or g8412 ( n16036 , n26178 , n437 );
    and g8413 ( n14297 , n11351 , n25765 );
    and g8414 ( n30030 , n26143 , n21001 );
    not g8415 ( n1328 , n20718 );
    not g8416 ( n13609 , n4571 );
    not g8417 ( n1983 , n479 );
    xnor g8418 ( n11999 , n22834 , n30650 );
    not g8419 ( n5452 , n15771 );
    xnor g8420 ( n20687 , n16883 , n21139 );
    or g8421 ( n47 , n26957 , n8757 );
    or g8422 ( n26417 , n31352 , n25591 );
    or g8423 ( n8548 , n25749 , n25399 );
    or g8424 ( n26211 , n2883 , n16177 );
    or g8425 ( n17022 , n1169 , n7569 );
    nor g8426 ( n4429 , n19366 , n19734 );
    or g8427 ( n4954 , n10340 , n23066 );
    xor g8428 ( n20676 , n23270 , n12566 );
    and g8429 ( n4725 , n16106 , n20986 );
    nor g8430 ( n10685 , n1039 , n2894 );
    or g8431 ( n17522 , n6036 , n27883 );
    not g8432 ( n15211 , n6063 );
    xnor g8433 ( n15829 , n16373 , n26392 );
    and g8434 ( n26820 , n16699 , n3470 );
    or g8435 ( n19447 , n31892 , n24934 );
    xnor g8436 ( n19594 , n4259 , n17945 );
    xor g8437 ( n30503 , n8575 , n5935 );
    or g8438 ( n1533 , n11262 , n22434 );
    or g8439 ( n16451 , n3268 , n15563 );
    and g8440 ( n31846 , n14193 , n21224 );
    or g8441 ( n21724 , n8293 , n11623 );
    or g8442 ( n7964 , n514 , n9448 );
    not g8443 ( n4457 , n3399 );
    and g8444 ( n7841 , n26864 , n29136 );
    buf g8445 ( n31070 , n26494 );
    xnor g8446 ( n31512 , n12208 , n14318 );
    xnor g8447 ( n31339 , n667 , n823 );
    xnor g8448 ( n24953 , n502 , n8407 );
    xnor g8449 ( n322 , n11079 , n31615 );
    or g8450 ( n19952 , n7955 , n22494 );
    and g8451 ( n6614 , n17948 , n15676 );
    and g8452 ( n31890 , n3135 , n18452 );
    not g8453 ( n22254 , n4238 );
    or g8454 ( n22482 , n7646 , n32 );
    xnor g8455 ( n11894 , n11241 , n12399 );
    or g8456 ( n9042 , n19024 , n8723 );
    not g8457 ( n10543 , n7124 );
    xnor g8458 ( n30074 , n9256 , n25020 );
    or g8459 ( n25312 , n1839 , n11120 );
    xnor g8460 ( n24080 , n24340 , n17438 );
    or g8461 ( n12469 , n22678 , n17411 );
    or g8462 ( n5185 , n29066 , n20740 );
    and g8463 ( n2895 , n16928 , n13359 );
    or g8464 ( n5565 , n13062 , n27881 );
    not g8465 ( n3711 , n1550 );
    xnor g8466 ( n28557 , n1975 , n7005 );
    xnor g8467 ( n18541 , n19752 , n22971 );
    or g8468 ( n31468 , n7184 , n9021 );
    or g8469 ( n16246 , n22023 , n23492 );
    not g8470 ( n18451 , n5813 );
    xnor g8471 ( n14161 , n19101 , n18388 );
    xnor g8472 ( n2159 , n29461 , n27342 );
    or g8473 ( n29729 , n280 , n30842 );
    or g8474 ( n28200 , n6712 , n8495 );
    xnor g8475 ( n5576 , n8974 , n23068 );
    xnor g8476 ( n23304 , n25568 , n18858 );
    xor g8477 ( n12508 , n9428 , n13434 );
    not g8478 ( n16987 , n26446 );
    and g8479 ( n15273 , n9448 , n514 );
    not g8480 ( n28327 , n23342 );
    not g8481 ( n19846 , n24503 );
    and g8482 ( n24071 , n26027 , n8976 );
    not g8483 ( n5322 , n8726 );
    or g8484 ( n9236 , n19624 , n19287 );
    and g8485 ( n24190 , n16377 , n31136 );
    not g8486 ( n15358 , n30633 );
    and g8487 ( n22432 , n25620 , n5880 );
    not g8488 ( n28108 , n26038 );
    and g8489 ( n18951 , n13505 , n2017 );
    not g8490 ( n8710 , n9894 );
    not g8491 ( n31389 , n3095 );
    not g8492 ( n4706 , n2623 );
    or g8493 ( n14057 , n724 , n27873 );
    not g8494 ( n9758 , n4978 );
    not g8495 ( n3459 , n13073 );
    or g8496 ( n24279 , n1281 , n16453 );
    or g8497 ( n28568 , n17508 , n18472 );
    or g8498 ( n20363 , n31555 , n20450 );
    not g8499 ( n31252 , n16111 );
    or g8500 ( n28785 , n17016 , n23638 );
    nor g8501 ( n19008 , n27292 , n23683 );
    or g8502 ( n28199 , n12446 , n20414 );
    or g8503 ( n16127 , n3643 , n6672 );
    xnor g8504 ( n29654 , n24856 , n16788 );
    not g8505 ( n14491 , n24258 );
    buf g8506 ( n29252 , n17233 );
    not g8507 ( n5090 , n27802 );
    or g8508 ( n11249 , n5948 , n8221 );
    xor g8509 ( n10398 , n22463 , n7529 );
    or g8510 ( n9641 , n21807 , n22003 );
    not g8511 ( n655 , n25889 );
    xnor g8512 ( n14569 , n21613 , n1692 );
    not g8513 ( n13597 , n9690 );
    xnor g8514 ( n24949 , n15675 , n18108 );
    xnor g8515 ( n14754 , n28551 , n18496 );
    and g8516 ( n26432 , n24082 , n5632 );
    not g8517 ( n2968 , n22242 );
    xnor g8518 ( n6694 , n10516 , n2973 );
    not g8519 ( n23508 , n19631 );
    xnor g8520 ( n3469 , n21745 , n29212 );
    xnor g8521 ( n14898 , n21617 , n24593 );
    xnor g8522 ( n2091 , n17824 , n21458 );
    not g8523 ( n142 , n22571 );
    not g8524 ( n10197 , n930 );
    not g8525 ( n9681 , n4226 );
    or g8526 ( n5972 , n27241 , n4497 );
    or g8527 ( n18321 , n1017 , n22860 );
    and g8528 ( n27680 , n7619 , n12625 );
    not g8529 ( n12743 , n15842 );
    not g8530 ( n7268 , n11826 );
    xnor g8531 ( n13222 , n1980 , n21808 );
    or g8532 ( n2254 , n14083 , n20093 );
    or g8533 ( n12590 , n24578 , n23585 );
    not g8534 ( n23640 , n22984 );
    xor g8535 ( n6963 , n11297 , n29945 );
    xnor g8536 ( n22641 , n7472 , n29684 );
    or g8537 ( n2807 , n4362 , n25867 );
    or g8538 ( n19932 , n23390 , n28693 );
    not g8539 ( n25004 , n25091 );
    xnor g8540 ( n4448 , n22841 , n1997 );
    xnor g8541 ( n12967 , n26029 , n256 );
    not g8542 ( n26414 , n7389 );
    not g8543 ( n28694 , n30090 );
    nor g8544 ( n1208 , n18832 , n31283 );
    xor g8545 ( n4487 , n23395 , n22431 );
    and g8546 ( n17925 , n9203 , n23072 );
    nor g8547 ( n23458 , n16986 , n27827 );
    and g8548 ( n7053 , n30499 , n26476 );
    nor g8549 ( n21557 , n7077 , n23646 );
    not g8550 ( n30099 , n11983 );
    xnor g8551 ( n16477 , n19220 , n19622 );
    nor g8552 ( n28215 , n26082 , n26445 );
    xnor g8553 ( n3816 , n19582 , n21960 );
    not g8554 ( n25069 , n9239 );
    or g8555 ( n27269 , n13436 , n19476 );
    and g8556 ( n25288 , n20603 , n3574 );
    and g8557 ( n24220 , n1989 , n598 );
    and g8558 ( n22779 , n23908 , n5048 );
    not g8559 ( n25704 , n17089 );
    or g8560 ( n4731 , n7013 , n11514 );
    xnor g8561 ( n31821 , n13466 , n31662 );
    xnor g8562 ( n6337 , n3355 , n10577 );
    and g8563 ( n22084 , n16473 , n8086 );
    nor g8564 ( n4152 , n25253 , n10776 );
    or g8565 ( n19527 , n31725 , n6429 );
    and g8566 ( n31523 , n7719 , n3876 );
    xnor g8567 ( n21234 , n10379 , n25152 );
    xnor g8568 ( n25424 , n21024 , n10570 );
    xor g8569 ( n17823 , n24208 , n15600 );
    nor g8570 ( n14813 , n23529 , n2591 );
    and g8571 ( n4097 , n16431 , n26754 );
    or g8572 ( n25420 , n14802 , n28063 );
    not g8573 ( n29966 , n23197 );
    and g8574 ( n15682 , n22663 , n24616 );
    not g8575 ( n5348 , n26308 );
    not g8576 ( n16773 , n28591 );
    not g8577 ( n6005 , n10142 );
    not g8578 ( n22279 , n167 );
    and g8579 ( n23460 , n6777 , n15536 );
    and g8580 ( n1972 , n12273 , n24444 );
    nor g8581 ( n26101 , n3149 , n9311 );
    xnor g8582 ( n906 , n29651 , n25657 );
    or g8583 ( n26837 , n9164 , n28294 );
    and g8584 ( n20652 , n11188 , n12952 );
    xor g8585 ( n24970 , n3929 , n13635 );
    xnor g8586 ( n1045 , n15065 , n22100 );
    or g8587 ( n7963 , n1282 , n2434 );
    xnor g8588 ( n7252 , n13330 , n13836 );
    not g8589 ( n8499 , n17866 );
    buf g8590 ( n11729 , n22367 );
    xor g8591 ( n9938 , n10396 , n4694 );
    or g8592 ( n26984 , n16467 , n26766 );
    or g8593 ( n17083 , n17617 , n11257 );
    xnor g8594 ( n23774 , n24209 , n9302 );
    and g8595 ( n28049 , n22312 , n2320 );
    xnor g8596 ( n1867 , n7450 , n22316 );
    not g8597 ( n23472 , n18072 );
    xnor g8598 ( n15756 , n28977 , n11267 );
    and g8599 ( n25964 , n24790 , n18386 );
    not g8600 ( n1204 , n6888 );
    nor g8601 ( n29165 , n30103 , n20344 );
    xnor g8602 ( n29257 , n19766 , n19359 );
    and g8603 ( n4440 , n2651 , n3431 );
    or g8604 ( n11081 , n5796 , n13890 );
    not g8605 ( n31327 , n1527 );
    xnor g8606 ( n3283 , n4741 , n3393 );
    and g8607 ( n19973 , n3903 , n30856 );
    xnor g8608 ( n12224 , n14939 , n20978 );
    not g8609 ( n25140 , n3492 );
    and g8610 ( n29326 , n2746 , n23171 );
    not g8611 ( n22835 , n30453 );
    xnor g8612 ( n13209 , n17131 , n5041 );
    or g8613 ( n25050 , n3635 , n22483 );
    nor g8614 ( n19130 , n20728 , n10259 );
    xnor g8615 ( n15190 , n21821 , n4703 );
    not g8616 ( n19879 , n21268 );
    and g8617 ( n4691 , n23863 , n23087 );
    and g8618 ( n9397 , n18476 , n18896 );
    not g8619 ( n24074 , n16678 );
    or g8620 ( n24538 , n27558 , n20738 );
    not g8621 ( n21292 , n2939 );
    and g8622 ( n26953 , n4670 , n25089 );
    nor g8623 ( n4841 , n21452 , n8846 );
    or g8624 ( n13199 , n1976 , n7689 );
    not g8625 ( n12211 , n14230 );
    nor g8626 ( n2854 , n14992 , n11197 );
    not g8627 ( n17645 , n19132 );
    or g8628 ( n10584 , n11796 , n1593 );
    not g8629 ( n26487 , n31007 );
    xnor g8630 ( n16728 , n24503 , n15396 );
    or g8631 ( n16808 , n23401 , n24584 );
    xnor g8632 ( n30575 , n23192 , n17821 );
    and g8633 ( n19744 , n31441 , n14478 );
    xnor g8634 ( n28821 , n5674 , n3745 );
    nor g8635 ( n6521 , n19392 , n24998 );
    and g8636 ( n21617 , n12964 , n21897 );
    nor g8637 ( n9255 , n22184 , n1886 );
    not g8638 ( n13054 , n2027 );
    xnor g8639 ( n1358 , n8488 , n23135 );
    and g8640 ( n8974 , n26030 , n8868 );
    not g8641 ( n11261 , n23131 );
    xor g8642 ( n30728 , n10648 , n30469 );
    or g8643 ( n18201 , n4245 , n13384 );
    or g8644 ( n24419 , n1146 , n20574 );
    and g8645 ( n25912 , n31971 , n9851 );
    not g8646 ( n25384 , n30817 );
    not g8647 ( n9097 , n3910 );
    not g8648 ( n2064 , n30366 );
    and g8649 ( n28148 , n3584 , n5717 );
    xnor g8650 ( n1411 , n31080 , n9729 );
    xnor g8651 ( n12188 , n9993 , n9723 );
    not g8652 ( n1190 , n9101 );
    and g8653 ( n24998 , n14143 , n6776 );
    or g8654 ( n6178 , n23709 , n12505 );
    not g8655 ( n14887 , n19299 );
    xnor g8656 ( n12767 , n22423 , n27591 );
    not g8657 ( n25203 , n20052 );
    xnor g8658 ( n24900 , n13367 , n30931 );
    xnor g8659 ( n3522 , n16083 , n7024 );
    xnor g8660 ( n31368 , n8154 , n8054 );
    not g8661 ( n14067 , n24827 );
    xor g8662 ( n8430 , n20709 , n28220 );
    or g8663 ( n22945 , n13343 , n11579 );
    not g8664 ( n19844 , n2991 );
    xnor g8665 ( n28958 , n8874 , n11051 );
    not g8666 ( n23574 , n6943 );
    xnor g8667 ( n9661 , n7705 , n31111 );
    or g8668 ( n30727 , n24702 , n14381 );
    and g8669 ( n29575 , n11104 , n25219 );
    xnor g8670 ( n16671 , n22768 , n29811 );
    or g8671 ( n12538 , n24757 , n5302 );
    xnor g8672 ( n22875 , n25929 , n26758 );
    not g8673 ( n11453 , n19196 );
    xnor g8674 ( n19746 , n25814 , n8407 );
    xnor g8675 ( n1809 , n28540 , n18981 );
    xnor g8676 ( n26343 , n28279 , n17462 );
    xnor g8677 ( n19424 , n25524 , n6928 );
    xnor g8678 ( n20570 , n8555 , n25984 );
    xnor g8679 ( n1279 , n12755 , n30239 );
    or g8680 ( n12491 , n10493 , n23982 );
    and g8681 ( n2773 , n6684 , n21917 );
    xnor g8682 ( n5701 , n18127 , n4214 );
    or g8683 ( n3061 , n16940 , n12793 );
    and g8684 ( n6455 , n9357 , n29519 );
    not g8685 ( n27008 , n6626 );
    or g8686 ( n5296 , n31722 , n28314 );
    xnor g8687 ( n10817 , n1920 , n4474 );
    xnor g8688 ( n29269 , n30464 , n6626 );
    xnor g8689 ( n21777 , n21112 , n4225 );
    xnor g8690 ( n22475 , n15588 , n24837 );
    or g8691 ( n23042 , n18534 , n25595 );
    xnor g8692 ( n26297 , n7705 , n10158 );
    xnor g8693 ( n31101 , n21623 , n23621 );
    not g8694 ( n4834 , n10802 );
    or g8695 ( n5764 , n11259 , n12230 );
    and g8696 ( n14987 , n10869 , n20975 );
    and g8697 ( n28649 , n8894 , n14444 );
    not g8698 ( n15255 , n8426 );
    or g8699 ( n29311 , n12002 , n28605 );
    or g8700 ( n22862 , n12783 , n8700 );
    not g8701 ( n26158 , n5101 );
    not g8702 ( n25569 , n22902 );
    and g8703 ( n30098 , n22629 , n8140 );
    and g8704 ( n24667 , n22689 , n13579 );
    xnor g8705 ( n31616 , n4283 , n30648 );
    not g8706 ( n11944 , n22537 );
    or g8707 ( n27197 , n13542 , n13628 );
    xnor g8708 ( n29607 , n15969 , n13786 );
    not g8709 ( n7575 , n16008 );
    and g8710 ( n16295 , n13292 , n31773 );
    not g8711 ( n6766 , n5902 );
    not g8712 ( n6238 , n4451 );
    or g8713 ( n9790 , n14916 , n30151 );
    or g8714 ( n15389 , n28113 , n14949 );
    xnor g8715 ( n16916 , n5395 , n23245 );
    or g8716 ( n5623 , n719 , n8980 );
    xor g8717 ( n13999 , n31106 , n14188 );
    not g8718 ( n11617 , n4344 );
    or g8719 ( n1684 , n27734 , n29496 );
    xnor g8720 ( n28067 , n30711 , n28807 );
    xnor g8721 ( n6224 , n27534 , n13725 );
    xnor g8722 ( n28739 , n13060 , n19315 );
    or g8723 ( n2260 , n17861 , n24572 );
    or g8724 ( n28547 , n18391 , n10952 );
    not g8725 ( n3395 , n30069 );
    and g8726 ( n7845 , n8735 , n10485 );
    and g8727 ( n23175 , n18822 , n4203 );
    xnor g8728 ( n21142 , n23678 , n27885 );
    or g8729 ( n6570 , n26629 , n13077 );
    xnor g8730 ( n10209 , n15225 , n14045 );
    and g8731 ( n14874 , n21173 , n3036 );
    xnor g8732 ( n21540 , n15347 , n20598 );
    nor g8733 ( n3298 , n6184 , n23818 );
    or g8734 ( n9647 , n3298 , n16615 );
    nor g8735 ( n16400 , n19935 , n965 );
    not g8736 ( n2450 , n27961 );
    not g8737 ( n559 , n19092 );
    or g8738 ( n20875 , n15249 , n27142 );
    or g8739 ( n13227 , n26942 , n13774 );
    or g8740 ( n1200 , n29987 , n4247 );
    xnor g8741 ( n8159 , n24881 , n6198 );
    and g8742 ( n26471 , n18666 , n9017 );
    not g8743 ( n963 , n27304 );
    nor g8744 ( n2980 , n8445 , n25883 );
    or g8745 ( n15900 , n15871 , n9872 );
    or g8746 ( n12171 , n2604 , n12162 );
    not g8747 ( n10730 , n1903 );
    not g8748 ( n6565 , n28674 );
    not g8749 ( n25239 , n20105 );
    not g8750 ( n10911 , n31002 );
    xnor g8751 ( n3793 , n24862 , n4774 );
    xnor g8752 ( n29859 , n12580 , n15669 );
    or g8753 ( n10098 , n31713 , n27648 );
    not g8754 ( n19322 , n21819 );
    nor g8755 ( n3378 , n20149 , n26756 );
    or g8756 ( n18162 , n19603 , n6262 );
    xnor g8757 ( n17968 , n29204 , n11887 );
    and g8758 ( n7126 , n12152 , n4548 );
    and g8759 ( n16037 , n10011 , n8227 );
    xor g8760 ( n21591 , n2679 , n28055 );
    and g8761 ( n19660 , n19267 , n29626 );
    not g8762 ( n14838 , n2686 );
    or g8763 ( n24506 , n16570 , n13167 );
    and g8764 ( n6559 , n343 , n29943 );
    or g8765 ( n30439 , n16411 , n3980 );
    or g8766 ( n29209 , n30584 , n19659 );
    and g8767 ( n25099 , n25599 , n8273 );
    not g8768 ( n18855 , n29084 );
    or g8769 ( n19327 , n24929 , n6038 );
    xnor g8770 ( n18204 , n26851 , n2916 );
    buf g8771 ( n6097 , n20364 );
    not g8772 ( n9882 , n101 );
    nor g8773 ( n20582 , n30961 , n946 );
    or g8774 ( n9584 , n14078 , n3776 );
    or g8775 ( n3421 , n31767 , n7721 );
    not g8776 ( n24613 , n13203 );
    or g8777 ( n18674 , n11918 , n25984 );
    not g8778 ( n4009 , n24304 );
    not g8779 ( n22396 , n18150 );
    not g8780 ( n18361 , n8681 );
    and g8781 ( n22618 , n9327 , n18059 );
    not g8782 ( n18668 , n26828 );
    and g8783 ( n1336 , n5874 , n25090 );
    xnor g8784 ( n6096 , n5638 , n11253 );
    xnor g8785 ( n25318 , n3801 , n20766 );
    xnor g8786 ( n5439 , n7314 , n31722 );
    nor g8787 ( n25010 , n26723 , n11798 );
    not g8788 ( n28262 , n20687 );
    xnor g8789 ( n18033 , n20785 , n1170 );
    or g8790 ( n25854 , n28810 , n24954 );
    xnor g8791 ( n21834 , n29390 , n24569 );
    or g8792 ( n3208 , n25491 , n28804 );
    xnor g8793 ( n15933 , n11360 , n9338 );
    or g8794 ( n10719 , n9941 , n29371 );
    xnor g8795 ( n8132 , n13307 , n29456 );
    nor g8796 ( n9052 , n26801 , n30376 );
    and g8797 ( n15090 , n6455 , n13476 );
    not g8798 ( n8878 , n12087 );
    not g8799 ( n25421 , n31679 );
    and g8800 ( n25796 , n29570 , n20736 );
    and g8801 ( n18232 , n11672 , n24578 );
    xnor g8802 ( n2429 , n6036 , n18207 );
    not g8803 ( n28825 , n31623 );
    or g8804 ( n11409 , n13582 , n27364 );
    nor g8805 ( n12553 , n11666 , n9565 );
    or g8806 ( n22705 , n15342 , n12860 );
    and g8807 ( n2362 , n3227 , n3538 );
    or g8808 ( n27624 , n27304 , n19288 );
    or g8809 ( n5464 , n15558 , n17878 );
    and g8810 ( n14997 , n18420 , n1691 );
    not g8811 ( n9967 , n23861 );
    not g8812 ( n23529 , n19808 );
    and g8813 ( n15277 , n24870 , n1392 );
    not g8814 ( n8255 , n29668 );
    and g8815 ( n16796 , n20355 , n17870 );
    and g8816 ( n8473 , n24905 , n18582 );
    or g8817 ( n26985 , n9939 , n8612 );
    or g8818 ( n11095 , n27233 , n22039 );
    not g8819 ( n29118 , n23716 );
    and g8820 ( n9335 , n22171 , n2581 );
    xnor g8821 ( n12564 , n2266 , n28558 );
    or g8822 ( n30440 , n7552 , n18731 );
    not g8823 ( n18403 , n24361 );
    not g8824 ( n30913 , n13555 );
    not g8825 ( n675 , n5873 );
    xnor g8826 ( n25413 , n11847 , n2825 );
    and g8827 ( n18876 , n30207 , n3765 );
    not g8828 ( n7220 , n24449 );
    nor g8829 ( n16279 , n14690 , n10269 );
    xnor g8830 ( n16196 , n24141 , n3059 );
    or g8831 ( n9950 , n7848 , n11888 );
    and g8832 ( n5889 , n31504 , n11095 );
    xnor g8833 ( n28589 , n8241 , n7664 );
    and g8834 ( n12492 , n12437 , n31338 );
    and g8835 ( n2374 , n18137 , n15395 );
    xnor g8836 ( n1745 , n18907 , n11866 );
    xnor g8837 ( n15400 , n22451 , n30908 );
    not g8838 ( n8509 , n29808 );
    xnor g8839 ( n30714 , n19142 , n27126 );
    and g8840 ( n5468 , n21189 , n24805 );
    nor g8841 ( n26944 , n22922 , n24066 );
    and g8842 ( n8832 , n31126 , n14772 );
    not g8843 ( n19029 , n6697 );
    xnor g8844 ( n21964 , n8092 , n9171 );
    nor g8845 ( n277 , n80 , n29874 );
    and g8846 ( n3472 , n5730 , n22241 );
    not g8847 ( n3123 , n6767 );
    xnor g8848 ( n13703 , n16337 , n1694 );
    not g8849 ( n23488 , n27613 );
    or g8850 ( n14632 , n6945 , n29731 );
    xnor g8851 ( n23835 , n18540 , n7475 );
    not g8852 ( n18940 , n19134 );
    or g8853 ( n7446 , n5156 , n20959 );
    or g8854 ( n25025 , n24727 , n16679 );
    nor g8855 ( n28335 , n26805 , n23911 );
    xor g8856 ( n21068 , n24653 , n26196 );
    nor g8857 ( n10440 , n15997 , n3311 );
    not g8858 ( n19245 , n12207 );
    and g8859 ( n24477 , n14074 , n12342 );
    not g8860 ( n166 , n7503 );
    xor g8861 ( n27492 , n7774 , n18003 );
    or g8862 ( n11534 , n14890 , n22313 );
    or g8863 ( n26588 , n28782 , n16056 );
    or g8864 ( n21398 , n18849 , n14701 );
    nor g8865 ( n19741 , n21544 , n2844 );
    not g8866 ( n23843 , n7482 );
    not g8867 ( n29188 , n9806 );
    xnor g8868 ( n18528 , n16045 , n20759 );
    and g8869 ( n23350 , n10538 , n2100 );
    or g8870 ( n7279 , n15999 , n9909 );
    and g8871 ( n11096 , n23106 , n7945 );
    nor g8872 ( n24309 , n12998 , n13410 );
    not g8873 ( n28136 , n19590 );
    or g8874 ( n9248 , n10076 , n29927 );
    or g8875 ( n5600 , n20784 , n22374 );
    xnor g8876 ( n21299 , n19265 , n10278 );
    xnor g8877 ( n8920 , n20057 , n21064 );
    xor g8878 ( n7574 , n11216 , n31723 );
    not g8879 ( n11666 , n30688 );
    not g8880 ( n9968 , n3166 );
    not g8881 ( n21585 , n12903 );
    xnor g8882 ( n16223 , n7734 , n15806 );
    and g8883 ( n16466 , n1374 , n16726 );
    not g8884 ( n14766 , n6642 );
    nor g8885 ( n9954 , n6180 , n28499 );
    and g8886 ( n23150 , n4857 , n31985 );
    and g8887 ( n30132 , n6257 , n3070 );
    nor g8888 ( n19226 , n1299 , n2334 );
    or g8889 ( n18226 , n18565 , n13675 );
    or g8890 ( n13492 , n24519 , n27598 );
    or g8891 ( n31011 , n13773 , n27863 );
    not g8892 ( n8638 , n8477 );
    or g8893 ( n12620 , n14484 , n16233 );
    nor g8894 ( n13753 , n15306 , n24275 );
    or g8895 ( n27669 , n19821 , n29340 );
    or g8896 ( n19578 , n15305 , n29824 );
    not g8897 ( n5599 , n4844 );
    not g8898 ( n12430 , n212 );
    not g8899 ( n14536 , n23520 );
    or g8900 ( n5245 , n7944 , n30447 );
    and g8901 ( n5397 , n31405 , n13369 );
    or g8902 ( n8382 , n16621 , n3673 );
    not g8903 ( n4591 , n19681 );
    xnor g8904 ( n2526 , n27647 , n6584 );
    not g8905 ( n11834 , n29367 );
    or g8906 ( n9570 , n4069 , n10879 );
    nor g8907 ( n2868 , n17841 , n10814 );
    xnor g8908 ( n5575 , n24445 , n21122 );
    nor g8909 ( n10605 , n15593 , n5567 );
    and g8910 ( n9636 , n26196 , n20486 );
    xnor g8911 ( n19533 , n31947 , n31206 );
    and g8912 ( n20896 , n11024 , n25107 );
    xnor g8913 ( n6836 , n28486 , n20430 );
    or g8914 ( n19272 , n26955 , n20174 );
    not g8915 ( n4469 , n10937 );
    xnor g8916 ( n28188 , n13455 , n24626 );
    or g8917 ( n31304 , n25879 , n13919 );
    xnor g8918 ( n11549 , n19071 , n18048 );
    not g8919 ( n28806 , n5241 );
    and g8920 ( n22953 , n23328 , n31877 );
    nor g8921 ( n5447 , n3735 , n17503 );
    xnor g8922 ( n6098 , n8911 , n29399 );
    nor g8923 ( n31700 , n8714 , n27919 );
    xnor g8924 ( n19334 , n15075 , n9604 );
    and g8925 ( n439 , n11559 , n27568 );
    xnor g8926 ( n892 , n554 , n5251 );
    or g8927 ( n31017 , n24026 , n14055 );
    and g8928 ( n171 , n23726 , n8030 );
    or g8929 ( n6323 , n21364 , n22481 );
    and g8930 ( n3826 , n25357 , n6215 );
    not g8931 ( n6315 , n21458 );
    nor g8932 ( n23709 , n12192 , n15095 );
    and g8933 ( n576 , n1959 , n22515 );
    xnor g8934 ( n3850 , n25175 , n5387 );
    and g8935 ( n23235 , n25200 , n30481 );
    and g8936 ( n18095 , n17746 , n29059 );
    and g8937 ( n13807 , n21543 , n20551 );
    or g8938 ( n8543 , n29975 , n4115 );
    not g8939 ( n12061 , n26798 );
    xnor g8940 ( n6659 , n24499 , n15983 );
    xnor g8941 ( n21028 , n17923 , n1923 );
    or g8942 ( n30157 , n15382 , n3171 );
    or g8943 ( n22364 , n24384 , n24542 );
    not g8944 ( n28795 , n22587 );
    or g8945 ( n26003 , n15949 , n18309 );
    or g8946 ( n3391 , n2620 , n14385 );
    not g8947 ( n25819 , n22807 );
    not g8948 ( n3572 , n9208 );
    xnor g8949 ( n22211 , n13462 , n19516 );
    or g8950 ( n24126 , n12625 , n944 );
    not g8951 ( n20923 , n16856 );
    or g8952 ( n82 , n25049 , n5696 );
    not g8953 ( n10200 , n5237 );
    not g8954 ( n12370 , n11223 );
    not g8955 ( n6411 , n28001 );
    not g8956 ( n12150 , n27088 );
    or g8957 ( n21147 , n23314 , n9184 );
    not g8958 ( n15235 , n10542 );
    and g8959 ( n17631 , n18717 , n26958 );
    and g8960 ( n4475 , n6723 , n22853 );
    nor g8961 ( n23305 , n1856 , n6633 );
    nor g8962 ( n19867 , n11373 , n31074 );
    not g8963 ( n3910 , n487 );
    not g8964 ( n14902 , n27301 );
    not g8965 ( n5578 , n20058 );
    xnor g8966 ( n25858 , n31247 , n21826 );
    xnor g8967 ( n5707 , n14040 , n561 );
    not g8968 ( n1327 , n31295 );
    nor g8969 ( n1129 , n1404 , n12533 );
    not g8970 ( n16710 , n8704 );
    xnor g8971 ( n19279 , n7985 , n27985 );
    and g8972 ( n8358 , n12042 , n31481 );
    not g8973 ( n10460 , n23453 );
    or g8974 ( n7370 , n5873 , n8087 );
    nor g8975 ( n14242 , n23556 , n14491 );
    not g8976 ( n28772 , n22836 );
    not g8977 ( n12630 , n8542 );
    not g8978 ( n8686 , n31094 );
    or g8979 ( n31008 , n12155 , n6814 );
    and g8980 ( n293 , n7973 , n10235 );
    and g8981 ( n3177 , n22359 , n9436 );
    xnor g8982 ( n2614 , n27421 , n5135 );
    or g8983 ( n21830 , n19953 , n1867 );
    or g8984 ( n20962 , n3191 , n727 );
    or g8985 ( n23988 , n22221 , n8488 );
    and g8986 ( n9747 , n27400 , n27480 );
    and g8987 ( n20290 , n17373 , n5606 );
    not g8988 ( n606 , n15342 );
    and g8989 ( n29354 , n8408 , n4772 );
    not g8990 ( n932 , n1084 );
    and g8991 ( n4963 , n18312 , n31019 );
    or g8992 ( n7700 , n4070 , n9769 );
    xnor g8993 ( n20989 , n5777 , n6925 );
    or g8994 ( n27773 , n1754 , n10016 );
    or g8995 ( n21148 , n6229 , n11212 );
    not g8996 ( n22210 , n16113 );
    or g8997 ( n14181 , n1347 , n20211 );
    xnor g8998 ( n21533 , n13993 , n29847 );
    and g8999 ( n16171 , n29171 , n19814 );
    not g9000 ( n25392 , n31982 );
    or g9001 ( n25341 , n10641 , n7256 );
    and g9002 ( n26509 , n16999 , n27269 );
    xnor g9003 ( n17430 , n26334 , n18399 );
    xnor g9004 ( n20631 , n22529 , n22294 );
    not g9005 ( n20439 , n14283 );
    not g9006 ( n14983 , n8496 );
    or g9007 ( n19968 , n29339 , n10698 );
    not g9008 ( n28217 , n4922 );
    xnor g9009 ( n29631 , n19103 , n31940 );
    not g9010 ( n29923 , n25272 );
    or g9011 ( n31581 , n6088 , n4636 );
    not g9012 ( n17197 , n13955 );
    and g9013 ( n5325 , n25181 , n2863 );
    xnor g9014 ( n6074 , n17129 , n11428 );
    xnor g9015 ( n4952 , n957 , n10101 );
    or g9016 ( n15832 , n9685 , n20207 );
    and g9017 ( n1780 , n17685 , n29605 );
    and g9018 ( n11004 , n14258 , n28995 );
    xnor g9019 ( n11477 , n31019 , n7760 );
    and g9020 ( n10588 , n7510 , n2903 );
    nor g9021 ( n806 , n6534 , n1831 );
    not g9022 ( n21057 , n793 );
    or g9023 ( n2208 , n19450 , n16823 );
    nor g9024 ( n16069 , n1856 , n11916 );
    and g9025 ( n16301 , n325 , n234 );
    xnor g9026 ( n15156 , n21944 , n7232 );
    and g9027 ( n19912 , n25611 , n5823 );
    xnor g9028 ( n29402 , n6187 , n9291 );
    not g9029 ( n6597 , n3782 );
    xnor g9030 ( n7675 , n29214 , n9675 );
    xnor g9031 ( n5521 , n25151 , n23118 );
    not g9032 ( n1082 , n14912 );
    xor g9033 ( n5962 , n4005 , n29807 );
    or g9034 ( n9081 , n31252 , n16375 );
    xnor g9035 ( n6971 , n26456 , n8042 );
    not g9036 ( n26277 , n9904 );
    xnor g9037 ( n30729 , n24982 , n4784 );
    and g9038 ( n20387 , n29572 , n20193 );
    xnor g9039 ( n15771 , n28184 , n12943 );
    and g9040 ( n15942 , n20932 , n1617 );
    and g9041 ( n2252 , n10757 , n25884 );
    not g9042 ( n13335 , n11507 );
    xnor g9043 ( n15842 , n29964 , n12478 );
    xnor g9044 ( n1475 , n29704 , n21758 );
    or g9045 ( n1332 , n11492 , n28931 );
    or g9046 ( n16049 , n29965 , n7138 );
    and g9047 ( n24572 , n7237 , n17534 );
    xnor g9048 ( n11733 , n9197 , n18419 );
    or g9049 ( n3231 , n24875 , n23684 );
    xor g9050 ( n20325 , n28430 , n16980 );
    xnor g9051 ( n1198 , n12675 , n116 );
    nor g9052 ( n16521 , n24638 , n8220 );
    not g9053 ( n14437 , n10269 );
    xnor g9054 ( n4199 , n10700 , n25011 );
    xnor g9055 ( n3680 , n27883 , n26002 );
    and g9056 ( n13917 , n1472 , n16504 );
    and g9057 ( n13228 , n15615 , n10834 );
    not g9058 ( n25165 , n2678 );
    and g9059 ( n3660 , n24052 , n12833 );
    and g9060 ( n23815 , n18353 , n20699 );
    and g9061 ( n23679 , n14517 , n17909 );
    or g9062 ( n11141 , n20521 , n20807 );
    nor g9063 ( n6088 , n554 , n23232 );
    or g9064 ( n6758 , n6181 , n12970 );
    xnor g9065 ( n15463 , n2528 , n24225 );
    or g9066 ( n2748 , n9491 , n28982 );
    not g9067 ( n22645 , n30163 );
    not g9068 ( n10219 , n31694 );
    or g9069 ( n22884 , n16177 , n12299 );
    or g9070 ( n2881 , n20926 , n18097 );
    or g9071 ( n8552 , n29356 , n30893 );
    nor g9072 ( n31606 , n6223 , n471 );
    xnor g9073 ( n8297 , n4191 , n7192 );
    xnor g9074 ( n9629 , n3438 , n1039 );
    or g9075 ( n25676 , n2653 , n5471 );
    or g9076 ( n18354 , n24309 , n1248 );
    xnor g9077 ( n7800 , n29059 , n27233 );
    not g9078 ( n24921 , n20567 );
    and g9079 ( n3992 , n7715 , n14432 );
    and g9080 ( n11952 , n21983 , n28785 );
    or g9081 ( n24259 , n1238 , n3410 );
    xnor g9082 ( n6549 , n23413 , n4673 );
    and g9083 ( n22002 , n13526 , n14227 );
    xor g9084 ( n28013 , n3945 , n19066 );
    and g9085 ( n8683 , n7748 , n17194 );
    xnor g9086 ( n943 , n5069 , n16815 );
    not g9087 ( n29590 , n19824 );
    xnor g9088 ( n1858 , n903 , n3008 );
    not g9089 ( n4143 , n18688 );
    xnor g9090 ( n21229 , n27105 , n30364 );
    not g9091 ( n17624 , n19386 );
    not g9092 ( n22149 , n405 );
    not g9093 ( n16413 , n20599 );
    xnor g9094 ( n29886 , n4970 , n16511 );
    nor g9095 ( n12666 , n24920 , n6750 );
    nor g9096 ( n23397 , n12983 , n28955 );
    and g9097 ( n25243 , n21972 , n15241 );
    or g9098 ( n16715 , n24404 , n19692 );
    or g9099 ( n5717 , n24753 , n30215 );
    xnor g9100 ( n21166 , n21199 , n8058 );
    not g9101 ( n27301 , n23949 );
    not g9102 ( n27661 , n24080 );
    not g9103 ( n12999 , n27186 );
    and g9104 ( n31939 , n28997 , n18021 );
    not g9105 ( n17803 , n20480 );
    xnor g9106 ( n18005 , n9744 , n11060 );
    and g9107 ( n31187 , n18969 , n19738 );
    and g9108 ( n4233 , n19065 , n27894 );
    xnor g9109 ( n22122 , n763 , n14361 );
    not g9110 ( n26904 , n19339 );
    not g9111 ( n18384 , n366 );
    xnor g9112 ( n21182 , n26147 , n2784 );
    and g9113 ( n13088 , n26046 , n10086 );
    xnor g9114 ( n12870 , n17292 , n29736 );
    nor g9115 ( n29989 , n29168 , n25324 );
    xnor g9116 ( n26920 , n24925 , n29361 );
    and g9117 ( n16899 , n20511 , n17701 );
    or g9118 ( n2083 , n3355 , n30971 );
    or g9119 ( n15513 , n27577 , n8789 );
    not g9120 ( n24439 , n19649 );
    and g9121 ( n444 , n10265 , n20769 );
    not g9122 ( n26826 , n14149 );
    not g9123 ( n15576 , n1315 );
    not g9124 ( n14149 , n8915 );
    not g9125 ( n30331 , n4286 );
    and g9126 ( n31195 , n13953 , n31449 );
    or g9127 ( n881 , n2539 , n22319 );
    nor g9128 ( n7923 , n26191 , n713 );
    not g9129 ( n11799 , n167 );
    and g9130 ( n9719 , n16990 , n2996 );
    xnor g9131 ( n30704 , n6127 , n8407 );
    or g9132 ( n4024 , n4170 , n18084 );
    and g9133 ( n15199 , n18268 , n7759 );
    or g9134 ( n4259 , n11136 , n31081 );
    nor g9135 ( n26244 , n29249 , n14480 );
    or g9136 ( n19486 , n521 , n29696 );
    nor g9137 ( n31805 , n11438 , n20604 );
    or g9138 ( n6519 , n1305 , n31097 );
    not g9139 ( n22059 , n23968 );
    and g9140 ( n4930 , n2806 , n22800 );
    not g9141 ( n20137 , n29157 );
    not g9142 ( n15362 , n14808 );
    not g9143 ( n28770 , n11866 );
    nor g9144 ( n5175 , n29390 , n24569 );
    or g9145 ( n23107 , n24638 , n7576 );
    not g9146 ( n3700 , n5809 );
    not g9147 ( n28857 , n16815 );
    or g9148 ( n2903 , n16724 , n28858 );
    buf g9149 ( n30865 , n30951 );
    or g9150 ( n10245 , n10735 , n20641 );
    and g9151 ( n1142 , n10256 , n5797 );
    not g9152 ( n13772 , n15737 );
    or g9153 ( n15160 , n31849 , n17405 );
    xnor g9154 ( n381 , n24512 , n24246 );
    not g9155 ( n28271 , n21182 );
    nor g9156 ( n5401 , n11601 , n28004 );
    nor g9157 ( n17191 , n1997 , n19493 );
    or g9158 ( n29505 , n6850 , n10145 );
    not g9159 ( n6481 , n9831 );
    xnor g9160 ( n27714 , n2464 , n15009 );
    xnor g9161 ( n11041 , n31725 , n11218 );
    or g9162 ( n13176 , n8407 , n23660 );
    nor g9163 ( n22760 , n25506 , n21258 );
    nor g9164 ( n14062 , n21846 , n27668 );
    or g9165 ( n16224 , n25545 , n24300 );
    or g9166 ( n18368 , n21458 , n30517 );
    or g9167 ( n4543 , n31436 , n19844 );
    or g9168 ( n6841 , n25089 , n12195 );
    xnor g9169 ( n2224 , n30562 , n20510 );
    or g9170 ( n11456 , n24525 , n11958 );
    or g9171 ( n7413 , n21960 , n28267 );
    not g9172 ( n9905 , n14595 );
    xnor g9173 ( n14548 , n14376 , n24246 );
    xnor g9174 ( n9494 , n30459 , n17981 );
    not g9175 ( n28800 , n11671 );
    xor g9176 ( n17141 , n20910 , n24036 );
    or g9177 ( n26214 , n27885 , n6209 );
    xnor g9178 ( n687 , n29755 , n246 );
    xor g9179 ( n19193 , n31501 , n8891 );
    not g9180 ( n10603 , n28268 );
    nor g9181 ( n21739 , n206 , n14061 );
    not g9182 ( n7520 , n31904 );
    not g9183 ( n21179 , n19667 );
    xnor g9184 ( n22601 , n13183 , n22369 );
    nor g9185 ( n20009 , n17910 , n7655 );
    xnor g9186 ( n1033 , n4181 , n12861 );
    not g9187 ( n19848 , n3281 );
    nor g9188 ( n21929 , n11368 , n14133 );
    not g9189 ( n14590 , n8079 );
    xnor g9190 ( n27566 , n16338 , n15892 );
    nor g9191 ( n27807 , n621 , n20190 );
    not g9192 ( n27820 , n24735 );
    xnor g9193 ( n9656 , n16167 , n27982 );
    and g9194 ( n18747 , n29221 , n13072 );
    or g9195 ( n13045 , n22422 , n30911 );
    not g9196 ( n7742 , n16367 );
    xnor g9197 ( n3546 , n28439 , n6110 );
    or g9198 ( n28446 , n23765 , n31096 );
    or g9199 ( n1041 , n17518 , n7472 );
    nor g9200 ( n9872 , n24664 , n25134 );
    not g9201 ( n19549 , n21749 );
    xnor g9202 ( n23431 , n28883 , n458 );
    or g9203 ( n31103 , n24055 , n19031 );
    xnor g9204 ( n4465 , n16404 , n16583 );
    nor g9205 ( n3093 , n19078 , n25346 );
    and g9206 ( n30048 , n2958 , n3086 );
    and g9207 ( n4839 , n2575 , n8648 );
    xnor g9208 ( n7092 , n20868 , n20330 );
    xnor g9209 ( n15550 , n23881 , n30672 );
    buf g9210 ( n7412 , n3906 );
    not g9211 ( n18555 , n25627 );
    not g9212 ( n9460 , n3062 );
    or g9213 ( n17701 , n21063 , n28624 );
    xnor g9214 ( n1752 , n28706 , n29144 );
    xnor g9215 ( n18042 , n31717 , n28161 );
    not g9216 ( n20999 , n16308 );
    and g9217 ( n5030 , n21696 , n14998 );
    or g9218 ( n7301 , n3798 , n31374 );
    and g9219 ( n9240 , n672 , n30706 );
    not g9220 ( n17021 , n17335 );
    not g9221 ( n196 , n10631 );
    or g9222 ( n26915 , n11341 , n15975 );
    and g9223 ( n2503 , n5587 , n29113 );
    nor g9224 ( n15337 , n6901 , n7052 );
    and g9225 ( n28248 , n15970 , n28231 );
    xnor g9226 ( n30640 , n30884 , n27737 );
    and g9227 ( n5724 , n14442 , n18049 );
    and g9228 ( n22840 , n27245 , n868 );
    not g9229 ( n17080 , n19094 );
    or g9230 ( n14652 , n7469 , n5391 );
    not g9231 ( n13478 , n12963 );
    not g9232 ( n8413 , n9202 );
    not g9233 ( n13875 , n11419 );
    nor g9234 ( n6282 , n14975 , n20572 );
    nor g9235 ( n510 , n6502 , n5208 );
    and g9236 ( n2929 , n28104 , n3741 );
    or g9237 ( n24737 , n17074 , n24517 );
    or g9238 ( n6762 , n29944 , n1978 );
    xnor g9239 ( n10084 , n15089 , n23441 );
    not g9240 ( n20717 , n27643 );
    or g9241 ( n7474 , n5016 , n24846 );
    or g9242 ( n21503 , n17232 , n29556 );
    or g9243 ( n6332 , n30514 , n15819 );
    buf g9244 ( n30651 , n25424 );
    not g9245 ( n29395 , n14076 );
    not g9246 ( n19449 , n23069 );
    not g9247 ( n27373 , n15121 );
    or g9248 ( n12835 , n29235 , n2833 );
    xnor g9249 ( n25272 , n6929 , n28691 );
    and g9250 ( n14524 , n22765 , n25063 );
    or g9251 ( n17891 , n16123 , n16759 );
    or g9252 ( n1492 , n10336 , n31437 );
    and g9253 ( n6319 , n5305 , n5069 );
    nor g9254 ( n29717 , n18955 , n7108 );
    and g9255 ( n10486 , n20835 , n28000 );
    not g9256 ( n18598 , n5836 );
    xnor g9257 ( n7037 , n29978 , n17019 );
    and g9258 ( n1290 , n30945 , n29141 );
    xnor g9259 ( n5221 , n3687 , n8043 );
    not g9260 ( n26641 , n28811 );
    or g9261 ( n27496 , n25677 , n4591 );
    not g9262 ( n30087 , n7082 );
    or g9263 ( n4356 , n28452 , n25394 );
    nor g9264 ( n19030 , n22149 , n6040 );
    not g9265 ( n23942 , n31653 );
    and g9266 ( n13573 , n25770 , n30885 );
    not g9267 ( n14441 , n27327 );
    or g9268 ( n10510 , n28482 , n2650 );
    and g9269 ( n14357 , n11176 , n10329 );
    and g9270 ( n12663 , n13927 , n16182 );
    xnor g9271 ( n4388 , n3650 , n5252 );
    not g9272 ( n17837 , n25291 );
    or g9273 ( n16490 , n4619 , n27026 );
    not g9274 ( n26449 , n18551 );
    or g9275 ( n12359 , n6911 , n21406 );
    or g9276 ( n28570 , n11092 , n24550 );
    xor g9277 ( n9088 , n11435 , n24687 );
    and g9278 ( n2136 , n19179 , n25334 );
    not g9279 ( n13463 , n28627 );
    or g9280 ( n12937 , n15739 , n5178 );
    nor g9281 ( n23944 , n23258 , n28463 );
    not g9282 ( n3724 , n29939 );
    and g9283 ( n20723 , n23249 , n23481 );
    not g9284 ( n29386 , n24879 );
    not g9285 ( n30601 , n7210 );
    nor g9286 ( n2826 , n2085 , n19581 );
    or g9287 ( n9272 , n1862 , n17683 );
    xnor g9288 ( n25018 , n17021 , n10593 );
    xnor g9289 ( n13444 , n2016 , n6719 );
    or g9290 ( n29700 , n28063 , n10312 );
    or g9291 ( n5005 , n11251 , n27268 );
    not g9292 ( n28003 , n24608 );
    and g9293 ( n10765 , n4413 , n15695 );
    or g9294 ( n22284 , n14411 , n17416 );
    xnor g9295 ( n22931 , n22922 , n19300 );
    or g9296 ( n11754 , n3213 , n27651 );
    or g9297 ( n19837 , n20481 , n16505 );
    or g9298 ( n31395 , n31222 , n18336 );
    buf g9299 ( n21137 , n20747 );
    not g9300 ( n25040 , n26294 );
    not g9301 ( n18836 , n8097 );
    nor g9302 ( n26125 , n23037 , n3197 );
    or g9303 ( n5145 , n6031 , n3060 );
    or g9304 ( n2941 , n23693 , n22019 );
    xnor g9305 ( n3913 , n16534 , n6750 );
    xnor g9306 ( n4569 , n17958 , n28626 );
    or g9307 ( n17436 , n10619 , n14861 );
    and g9308 ( n7116 , n22179 , n22686 );
    not g9309 ( n31049 , n1279 );
    buf g9310 ( n20067 , n4935 );
    not g9311 ( n10119 , n10881 );
    not g9312 ( n20360 , n11630 );
    or g9313 ( n8659 , n1046 , n17566 );
    xnor g9314 ( n19569 , n15440 , n22527 );
    xnor g9315 ( n21444 , n27822 , n1827 );
    xnor g9316 ( n9197 , n2380 , n8596 );
    and g9317 ( n15607 , n30200 , n28398 );
    or g9318 ( n9667 , n17661 , n6890 );
    nor g9319 ( n3887 , n17745 , n24068 );
    not g9320 ( n13201 , n12217 );
    or g9321 ( n23434 , n270 , n6051 );
    not g9322 ( n3295 , n27896 );
    and g9323 ( n5704 , n20335 , n6223 );
    and g9324 ( n26352 , n20556 , n460 );
    or g9325 ( n15086 , n28180 , n24002 );
    or g9326 ( n16704 , n24193 , n16316 );
    xnor g9327 ( n25718 , n2492 , n25267 );
    nor g9328 ( n28299 , n30255 , n21719 );
    and g9329 ( n685 , n10622 , n29726 );
    or g9330 ( n18787 , n7414 , n28697 );
    nor g9331 ( n6954 , n1863 , n12119 );
    xnor g9332 ( n2163 , n20186 , n18647 );
    and g9333 ( n20007 , n26851 , n18994 );
    not g9334 ( n25550 , n18246 );
    xnor g9335 ( n31263 , n18191 , n30115 );
    and g9336 ( n12070 , n11742 , n17692 );
    not g9337 ( n9342 , n25350 );
    not g9338 ( n12594 , n830 );
    not g9339 ( n19077 , n17341 );
    not g9340 ( n11340 , n22688 );
    xnor g9341 ( n30394 , n7136 , n14580 );
    or g9342 ( n5735 , n21162 , n23128 );
    or g9343 ( n19423 , n7317 , n19349 );
    not g9344 ( n20069 , n22731 );
    not g9345 ( n19733 , n17622 );
    nor g9346 ( n27711 , n17745 , n12920 );
    xnor g9347 ( n22666 , n25928 , n29976 );
    nor g9348 ( n12343 , n20601 , n16862 );
    nor g9349 ( n30240 , n27355 , n2116 );
    or g9350 ( n28941 , n25804 , n636 );
    and g9351 ( n6580 , n1470 , n22225 );
    not g9352 ( n20607 , n2802 );
    or g9353 ( n2822 , n19753 , n29214 );
    not g9354 ( n25183 , n23002 );
    not g9355 ( n21750 , n821 );
    or g9356 ( n1156 , n22831 , n24818 );
    or g9357 ( n26120 , n12998 , n2571 );
    not g9358 ( n31586 , n17089 );
    and g9359 ( n18760 , n24667 , n10423 );
    not g9360 ( n5938 , n29870 );
    not g9361 ( n9172 , n7928 );
    not g9362 ( n7995 , n5973 );
    xnor g9363 ( n21971 , n21631 , n31821 );
    or g9364 ( n29486 , n18197 , n10907 );
    xnor g9365 ( n23716 , n310 , n1064 );
    xnor g9366 ( n27556 , n14481 , n29564 );
    or g9367 ( n15621 , n22818 , n12820 );
    and g9368 ( n14511 , n28570 , n28383 );
    and g9369 ( n7329 , n19774 , n12662 );
    or g9370 ( n18625 , n30219 , n912 );
    or g9371 ( n14578 , n2312 , n30420 );
    not g9372 ( n25701 , n22088 );
    or g9373 ( n8375 , n8064 , n16977 );
    nor g9374 ( n22699 , n26004 , n10863 );
    not g9375 ( n14656 , n27708 );
    not g9376 ( n22398 , n8469 );
    xnor g9377 ( n5613 , n28910 , n3839 );
    not g9378 ( n8993 , n27774 );
    xnor g9379 ( n21372 , n15851 , n389 );
    or g9380 ( n13809 , n31317 , n11965 );
    and g9381 ( n29753 , n3100 , n25122 );
    nor g9382 ( n19061 , n15127 , n11850 );
    xnor g9383 ( n4408 , n17678 , n19587 );
    or g9384 ( n24267 , n19362 , n23664 );
    or g9385 ( n18874 , n16856 , n3265 );
    or g9386 ( n12162 , n964 , n407 );
    nor g9387 ( n7565 , n4711 , n9150 );
    not g9388 ( n26774 , n17682 );
    not g9389 ( n14289 , n6803 );
    xnor g9390 ( n6286 , n17979 , n14370 );
    or g9391 ( n11647 , n22286 , n24007 );
    and g9392 ( n10831 , n25051 , n29199 );
    not g9393 ( n13743 , n14426 );
    nor g9394 ( n12423 , n14690 , n26259 );
    and g9395 ( n3998 , n23169 , n15396 );
    not g9396 ( n3602 , n30336 );
    and g9397 ( n16903 , n30839 , n23049 );
    or g9398 ( n22155 , n4006 , n31412 );
    xnor g9399 ( n13763 , n4480 , n6957 );
    and g9400 ( n30781 , n8327 , n4607 );
    or g9401 ( n8859 , n6569 , n9289 );
    or g9402 ( n25019 , n6163 , n18257 );
    or g9403 ( n17017 , n30936 , n21814 );
    or g9404 ( n26064 , n2588 , n28114 );
    xnor g9405 ( n4626 , n26409 , n30568 );
    xor g9406 ( n12572 , n28853 , n5981 );
    not g9407 ( n28990 , n3747 );
    xnor g9408 ( n6890 , n9811 , n20159 );
    not g9409 ( n10637 , n29849 );
    xnor g9410 ( n31190 , n6367 , n31334 );
    and g9411 ( n3924 , n28945 , n5715 );
    buf g9412 ( n6560 , n28298 );
    and g9413 ( n21449 , n15442 , n26035 );
    xnor g9414 ( n20092 , n20791 , n8360 );
    and g9415 ( n11073 , n7557 , n10873 );
    or g9416 ( n2582 , n15185 , n12480 );
    or g9417 ( n8181 , n26240 , n17486 );
    and g9418 ( n9951 , n19163 , n26167 );
    and g9419 ( n2211 , n19287 , n21084 );
    buf g9420 ( n29368 , n2205 );
    xnor g9421 ( n17418 , n8457 , n8714 );
    nor g9422 ( n10609 , n3782 , n21308 );
    xnor g9423 ( n23987 , n6127 , n5948 );
    or g9424 ( n11398 , n8275 , n27418 );
    and g9425 ( n27376 , n28905 , n1936 );
    or g9426 ( n25489 , n2883 , n23727 );
    not g9427 ( n18596 , n12441 );
    or g9428 ( n22593 , n25458 , n19152 );
    and g9429 ( n26567 , n16247 , n25341 );
    or g9430 ( n27797 , n1518 , n6153 );
    nor g9431 ( n27094 , n21208 , n8907 );
    not g9432 ( n3655 , n4257 );
    not g9433 ( n15610 , n23927 );
    or g9434 ( n29997 , n10139 , n107 );
    nor g9435 ( n28961 , n27233 , n10751 );
    or g9436 ( n7523 , n29954 , n25602 );
    xor g9437 ( n28887 , n1705 , n18200 );
    or g9438 ( n31609 , n3883 , n5287 );
    not g9439 ( n9235 , n18389 );
    and g9440 ( n49 , n16850 , n11518 );
    or g9441 ( n5987 , n17019 , n6426 );
    and g9442 ( n2247 , n13805 , n11444 );
    xnor g9443 ( n21835 , n5743 , n11829 );
    not g9444 ( n8233 , n18840 );
    xnor g9445 ( n25825 , n31481 , n13859 );
    and g9446 ( n29508 , n5859 , n11107 );
    or g9447 ( n24950 , n14342 , n12353 );
    and g9448 ( n10361 , n21559 , n21652 );
    not g9449 ( n19004 , n18918 );
    not g9450 ( n2236 , n998 );
    not g9451 ( n17574 , n3606 );
    xnor g9452 ( n17086 , n12808 , n19118 );
    or g9453 ( n25732 , n8584 , n30828 );
    xnor g9454 ( n21844 , n4610 , n16079 );
    not g9455 ( n813 , n21063 );
    not g9456 ( n16294 , n3808 );
    and g9457 ( n16373 , n15385 , n30665 );
    xnor g9458 ( n26732 , n23789 , n26884 );
    or g9459 ( n9104 , n31501 , n7924 );
    or g9460 ( n9536 , n20222 , n23790 );
    not g9461 ( n13103 , n18366 );
    not g9462 ( n15962 , n2648 );
    xnor g9463 ( n28029 , n16096 , n1923 );
    and g9464 ( n13216 , n23583 , n12785 );
    not g9465 ( n11362 , n19434 );
    xnor g9466 ( n14163 , n19505 , n22142 );
    not g9467 ( n24514 , n16776 );
    xnor g9468 ( n23630 , n4524 , n31502 );
    and g9469 ( n11723 , n20865 , n6900 );
    xnor g9470 ( n4622 , n30299 , n30119 );
    or g9471 ( n12161 , n14736 , n28192 );
    and g9472 ( n7071 , n23710 , n15233 );
    and g9473 ( n4343 , n23953 , n17907 );
    and g9474 ( n27674 , n23708 , n18465 );
    or g9475 ( n2581 , n14950 , n7624 );
    and g9476 ( n193 , n30115 , n18191 );
    nor g9477 ( n30371 , n11239 , n14307 );
    xnor g9478 ( n8906 , n6767 , n2515 );
    xnor g9479 ( n22569 , n6221 , n17981 );
    not g9480 ( n24750 , n15698 );
    and g9481 ( n27583 , n15629 , n1643 );
    xnor g9482 ( n19995 , n7292 , n2536 );
    nor g9483 ( n22144 , n11886 , n1913 );
    or g9484 ( n31602 , n2227 , n13185 );
    xnor g9485 ( n31744 , n19900 , n10951 );
    not g9486 ( n26529 , n13210 );
    xor g9487 ( n3980 , n29979 , n5707 );
    xnor g9488 ( n22036 , n18915 , n8705 );
    not g9489 ( n1191 , n10468 );
    not g9490 ( n28280 , n29660 );
    xnor g9491 ( n27058 , n26784 , n22597 );
    xnor g9492 ( n17941 , n17214 , n19901 );
    not g9493 ( n21549 , n7262 );
    not g9494 ( n14736 , n18027 );
    not g9495 ( n29647 , n21488 );
    nor g9496 ( n18034 , n24990 , n22561 );
    or g9497 ( n22473 , n21667 , n20313 );
    or g9498 ( n768 , n20293 , n8446 );
    xnor g9499 ( n18851 , n17294 , n17046 );
    and g9500 ( n21128 , n18276 , n14673 );
    not g9501 ( n28535 , n23394 );
    and g9502 ( n20161 , n2819 , n15297 );
    or g9503 ( n27421 , n15087 , n2193 );
    and g9504 ( n4284 , n24409 , n25981 );
    or g9505 ( n19480 , n6176 , n31984 );
    not g9506 ( n15233 , n28638 );
    not g9507 ( n13398 , n12712 );
    or g9508 ( n11683 , n7055 , n14499 );
    nor g9509 ( n11793 , n21508 , n22981 );
    and g9510 ( n26465 , n4044 , n18674 );
    xnor g9511 ( n26668 , n26889 , n3272 );
    or g9512 ( n12336 , n9404 , n21450 );
    or g9513 ( n16939 , n24013 , n25159 );
    xnor g9514 ( n28898 , n11368 , n11601 );
    xnor g9515 ( n22729 , n23622 , n9879 );
    xnor g9516 ( n12455 , n11799 , n6349 );
    not g9517 ( n30681 , n13758 );
    nor g9518 ( n128 , n2794 , n8386 );
    and g9519 ( n1766 , n5171 , n21858 );
    xnor g9520 ( n20316 , n31204 , n30405 );
    xnor g9521 ( n5914 , n22832 , n23061 );
    or g9522 ( n7045 , n27069 , n11523 );
    nor g9523 ( n18325 , n15178 , n20922 );
    and g9524 ( n577 , n31554 , n16985 );
    xnor g9525 ( n11724 , n27544 , n21816 );
    not g9526 ( n7262 , n26623 );
    xnor g9527 ( n24010 , n27865 , n8561 );
    xnor g9528 ( n1376 , n20023 , n16767 );
    or g9529 ( n15522 , n25149 , n8545 );
    xnor g9530 ( n25786 , n28030 , n20483 );
    not g9531 ( n16296 , n22518 );
    or g9532 ( n4008 , n29264 , n281 );
    or g9533 ( n10613 , n24587 , n838 );
    xnor g9534 ( n12340 , n24685 , n13966 );
    or g9535 ( n21500 , n5715 , n28945 );
    not g9536 ( n7535 , n27534 );
    xnor g9537 ( n7155 , n24778 , n25331 );
    buf g9538 ( n4372 , n26771 );
    and g9539 ( n15587 , n21353 , n3707 );
    or g9540 ( n31236 , n1833 , n8015 );
    not g9541 ( n24332 , n30801 );
    or g9542 ( n20265 , n19381 , n7920 );
    xnor g9543 ( n1388 , n30140 , n9092 );
    xnor g9544 ( n9138 , n29199 , n24401 );
    not g9545 ( n29946 , n311 );
    or g9546 ( n18615 , n22347 , n19975 );
    or g9547 ( n31117 , n12343 , n7873 );
    and g9548 ( n8420 , n45 , n21031 );
    nor g9549 ( n14084 , n8321 , n28314 );
    xnor g9550 ( n15318 , n19197 , n2709 );
    xnor g9551 ( n29666 , n3852 , n23689 );
    not g9552 ( n23366 , n30976 );
    or g9553 ( n10771 , n1692 , n23666 );
    not g9554 ( n13414 , n2476 );
    not g9555 ( n25503 , n14777 );
    and g9556 ( n20956 , n14839 , n14534 );
    or g9557 ( n21222 , n10853 , n10713 );
    nor g9558 ( n3559 , n26390 , n11560 );
    xor g9559 ( n8301 , n3805 , n11860 );
    not g9560 ( n13973 , n1105 );
    xor g9561 ( n20545 , n4151 , n13512 );
    and g9562 ( n16964 , n16750 , n11683 );
    not g9563 ( n22800 , n25512 );
    not g9564 ( n14000 , n1130 );
    and g9565 ( n21382 , n1593 , n30099 );
    or g9566 ( n7786 , n12526 , n20216 );
    not g9567 ( n23418 , n26168 );
    nor g9568 ( n24521 , n8338 , n27918 );
    xnor g9569 ( n30772 , n5889 , n21073 );
    xnor g9570 ( n24244 , n19108 , n19631 );
    not g9571 ( n14965 , n19529 );
    not g9572 ( n21284 , n573 );
    or g9573 ( n22684 , n25906 , n8785 );
    not g9574 ( n25749 , n16283 );
    or g9575 ( n623 , n16855 , n31807 );
    or g9576 ( n24393 , n26652 , n18784 );
    and g9577 ( n2735 , n30559 , n20263 );
    or g9578 ( n11878 , n5412 , n31334 );
    xnor g9579 ( n7243 , n7651 , n14992 );
    not g9580 ( n22324 , n27176 );
    xnor g9581 ( n29276 , n11705 , n7651 );
    nor g9582 ( n18968 , n24525 , n19046 );
    not g9583 ( n9174 , n673 );
    xnor g9584 ( n30174 , n12321 , n11333 );
    nor g9585 ( n20621 , n15219 , n30102 );
    not g9586 ( n13680 , n20236 );
    xnor g9587 ( n23776 , n23616 , n7694 );
    and g9588 ( n31082 , n25241 , n19946 );
    xnor g9589 ( n8628 , n27312 , n15499 );
    not g9590 ( n14276 , n4911 );
    nor g9591 ( n27857 , n2759 , n5708 );
    nor g9592 ( n6400 , n8340 , n10277 );
    xnor g9593 ( n22836 , n1666 , n24010 );
    or g9594 ( n22584 , n4812 , n5556 );
    xnor g9595 ( n12165 , n12600 , n19323 );
    and g9596 ( n21168 , n15154 , n3530 );
    xnor g9597 ( n30792 , n11417 , n27471 );
    and g9598 ( n2761 , n11961 , n28696 );
    xnor g9599 ( n12253 , n30693 , n23799 );
    not g9600 ( n6450 , n18117 );
    not g9601 ( n9048 , n8032 );
    xnor g9602 ( n29186 , n19216 , n31883 );
    and g9603 ( n10007 , n3825 , n15355 );
    and g9604 ( n6328 , n23564 , n7911 );
    or g9605 ( n2837 , n31851 , n31274 );
    xnor g9606 ( n116 , n21069 , n329 );
    xor g9607 ( n6139 , n24256 , n28054 );
    xnor g9608 ( n14337 , n29402 , n14100 );
    xnor g9609 ( n13383 , n19293 , n13141 );
    or g9610 ( n10545 , n183 , n14019 );
    and g9611 ( n20285 , n15810 , n20208 );
    nor g9612 ( n14483 , n16812 , n13097 );
    and g9613 ( n14760 , n13652 , n26813 );
    xnor g9614 ( n474 , n2901 , n8223 );
    not g9615 ( n16086 , n17632 );
    or g9616 ( n26702 , n9515 , n16892 );
    or g9617 ( n14528 , n496 , n8880 );
    not g9618 ( n28026 , n14340 );
    and g9619 ( n11688 , n19643 , n8834 );
    or g9620 ( n6776 , n23725 , n13568 );
    xor g9621 ( n20473 , n798 , n5266 );
    nor g9622 ( n8279 , n12030 , n13378 );
    not g9623 ( n25745 , n2001 );
    xnor g9624 ( n16093 , n10700 , n7432 );
    and g9625 ( n30809 , n21691 , n25840 );
    xnor g9626 ( n6423 , n26761 , n31166 );
    and g9627 ( n625 , n27903 , n2465 );
    and g9628 ( n31808 , n13599 , n18960 );
    not g9629 ( n17346 , n7149 );
    not g9630 ( n17151 , n13120 );
    or g9631 ( n24688 , n25710 , n25511 );
    not g9632 ( n6681 , n24455 );
    and g9633 ( n2787 , n24203 , n31892 );
    not g9634 ( n10635 , n31524 );
    not g9635 ( n26359 , n1742 );
    and g9636 ( n29977 , n23794 , n2587 );
    and g9637 ( n8557 , n877 , n27333 );
    not g9638 ( n11295 , n26720 );
    xnor g9639 ( n5555 , n24574 , n11850 );
    xnor g9640 ( n28569 , n27902 , n3249 );
    or g9641 ( n6451 , n11317 , n24385 );
    or g9642 ( n13581 , n2629 , n6552 );
    or g9643 ( n4656 , n20453 , n19699 );
    not g9644 ( n10260 , n13331 );
    or g9645 ( n15850 , n22510 , n28296 );
    xnor g9646 ( n24739 , n29915 , n7809 );
    nor g9647 ( n6439 , n5361 , n19464 );
    xnor g9648 ( n22148 , n11658 , n16609 );
    or g9649 ( n30224 , n28327 , n18216 );
    xnor g9650 ( n66 , n9002 , n6370 );
    or g9651 ( n24282 , n4707 , n10717 );
    xnor g9652 ( n14593 , n22899 , n452 );
    or g9653 ( n22329 , n14150 , n12506 );
    xnor g9654 ( n3831 , n7879 , n19406 );
    not g9655 ( n22335 , n31170 );
    buf g9656 ( n28058 , n20020 );
    or g9657 ( n7601 , n23339 , n9138 );
    nor g9658 ( n4681 , n3205 , n28663 );
    not g9659 ( n12402 , n23813 );
    or g9660 ( n9506 , n15431 , n7566 );
    xnor g9661 ( n8298 , n30445 , n12181 );
    or g9662 ( n25645 , n6995 , n27205 );
    and g9663 ( n26788 , n14623 , n12703 );
    and g9664 ( n545 , n12241 , n13301 );
    not g9665 ( n29708 , n16604 );
    not g9666 ( n31634 , n24120 );
    not g9667 ( n26869 , n13429 );
    nor g9668 ( n17260 , n23077 , n21128 );
    or g9669 ( n29724 , n22012 , n25158 );
    or g9670 ( n15661 , n22010 , n18928 );
    xnor g9671 ( n2538 , n23910 , n1614 );
    and g9672 ( n15703 , n10418 , n18806 );
    nor g9673 ( n9875 , n12642 , n30085 );
    buf g9674 ( n27948 , n2858 );
    or g9675 ( n28130 , n25962 , n10010 );
    nor g9676 ( n8607 , n25760 , n16865 );
    xnor g9677 ( n9762 , n3907 , n15436 );
    nor g9678 ( n19415 , n18146 , n533 );
    or g9679 ( n1134 , n20978 , n30054 );
    or g9680 ( n16141 , n16829 , n23235 );
    not g9681 ( n25937 , n5332 );
    xnor g9682 ( n17492 , n368 , n8822 );
    or g9683 ( n8002 , n31722 , n14089 );
    or g9684 ( n2860 , n28365 , n13900 );
    not g9685 ( n28398 , n12673 );
    and g9686 ( n26356 , n3235 , n23379 );
    nor g9687 ( n5200 , n8017 , n26264 );
    xnor g9688 ( n19109 , n20200 , n344 );
    xnor g9689 ( n25946 , n2223 , n12936 );
    not g9690 ( n27650 , n6367 );
    xnor g9691 ( n27880 , n8620 , n29902 );
    nor g9692 ( n15533 , n28006 , n2511 );
    or g9693 ( n2737 , n21947 , n2072 );
    xnor g9694 ( n26660 , n29796 , n22233 );
    and g9695 ( n11977 , n3088 , n14384 );
    xnor g9696 ( n28640 , n6836 , n5559 );
    or g9697 ( n12648 , n6373 , n9897 );
    or g9698 ( n27903 , n3441 , n8215 );
    and g9699 ( n4319 , n23086 , n27059 );
    or g9700 ( n6932 , n30265 , n29161 );
    nor g9701 ( n29038 , n10071 , n20825 );
    xnor g9702 ( n6445 , n23721 , n12767 );
    and g9703 ( n31832 , n20695 , n24739 );
    xnor g9704 ( n6492 , n20951 , n17472 );
    xnor g9705 ( n29140 , n10264 , n21272 );
    xnor g9706 ( n13161 , n10265 , n6480 );
    nor g9707 ( n6853 , n15649 , n22811 );
    xnor g9708 ( n28259 , n17951 , n13121 );
    xnor g9709 ( n9026 , n27251 , n8901 );
    nor g9710 ( n2230 , n26082 , n6957 );
    buf g9711 ( n18259 , n26751 );
    or g9712 ( n14687 , n10327 , n8944 );
    and g9713 ( n27641 , n10850 , n1369 );
    or g9714 ( n29530 , n4662 , n7489 );
    or g9715 ( n18196 , n24631 , n27014 );
    xnor g9716 ( n24022 , n25431 , n8694 );
    not g9717 ( n26690 , n10348 );
    nor g9718 ( n28219 , n3641 , n31401 );
    xnor g9719 ( n12431 , n13957 , n15987 );
    not g9720 ( n20240 , n3338 );
    and g9721 ( n29712 , n16578 , n26049 );
    xnor g9722 ( n22708 , n23940 , n29846 );
    not g9723 ( n29961 , n13152 );
    not g9724 ( n30523 , n16096 );
    xor g9725 ( n2454 , n3582 , n30710 );
    not g9726 ( n28264 , n29444 );
    and g9727 ( n20411 , n11097 , n6792 );
    xnor g9728 ( n2004 , n12598 , n13029 );
    xnor g9729 ( n10932 , n29629 , n12392 );
    or g9730 ( n20506 , n21597 , n31435 );
    or g9731 ( n31985 , n10043 , n23591 );
    xnor g9732 ( n22405 , n22150 , n27959 );
    and g9733 ( n24498 , n9025 , n5541 );
    not g9734 ( n10187 , n16350 );
    xnor g9735 ( n2359 , n11615 , n12562 );
    or g9736 ( n17709 , n1991 , n9951 );
    or g9737 ( n4781 , n13287 , n17166 );
    or g9738 ( n29765 , n9163 , n25727 );
    or g9739 ( n29139 , n30411 , n17880 );
    or g9740 ( n6582 , n31737 , n3672 );
    and g9741 ( n7460 , n10752 , n18182 );
    xnor g9742 ( n8330 , n6447 , n20933 );
    not g9743 ( n18124 , n1794 );
    or g9744 ( n7088 , n267 , n1651 );
    or g9745 ( n19903 , n15930 , n30741 );
    nor g9746 ( n29738 , n25733 , n6521 );
    xnor g9747 ( n5089 , n11830 , n26906 );
    not g9748 ( n29965 , n23914 );
    xnor g9749 ( n17117 , n11971 , n7330 );
    and g9750 ( n31977 , n25631 , n28722 );
    not g9751 ( n18048 , n20364 );
    xnor g9752 ( n24724 , n30147 , n29514 );
    or g9753 ( n26958 , n13494 , n23897 );
    nor g9754 ( n10199 , n31718 , n16096 );
    or g9755 ( n23137 , n10645 , n28725 );
    xnor g9756 ( n13758 , n12667 , n4465 );
    and g9757 ( n7312 , n18888 , n8636 );
    xnor g9758 ( n12745 , n1774 , n3570 );
    or g9759 ( n1729 , n13974 , n10452 );
    xnor g9760 ( n27608 , n3097 , n28287 );
    xor g9761 ( n25596 , n22682 , n6258 );
    nor g9762 ( n17873 , n7656 , n12728 );
    and g9763 ( n10548 , n23056 , n21485 );
    not g9764 ( n11624 , n13957 );
    and g9765 ( n2725 , n24314 , n18628 );
    not g9766 ( n7947 , n6495 );
    and g9767 ( n30178 , n3980 , n16411 );
    or g9768 ( n27189 , n14997 , n13807 );
    or g9769 ( n5636 , n18289 , n13373 );
    xnor g9770 ( n5462 , n13229 , n19270 );
    not g9771 ( n31710 , n20717 );
    not g9772 ( n11635 , n11655 );
    or g9773 ( n27803 , n28523 , n5065 );
    not g9774 ( n20107 , n29432 );
    nor g9775 ( n13745 , n17995 , n1132 );
    xnor g9776 ( n17413 , n5582 , n27896 );
    or g9777 ( n24912 , n26191 , n18147 );
    or g9778 ( n23645 , n11216 , n22410 );
    not g9779 ( n25338 , n515 );
    and g9780 ( n17349 , n31225 , n24296 );
    not g9781 ( n21926 , n3641 );
    and g9782 ( n26835 , n19635 , n5070 );
    nor g9783 ( n2414 , n29897 , n7663 );
    xnor g9784 ( n11682 , n27726 , n8414 );
    not g9785 ( n10930 , n23861 );
    or g9786 ( n15637 , n8009 , n13132 );
    not g9787 ( n8573 , n23475 );
    or g9788 ( n26962 , n29820 , n31943 );
    not g9789 ( n1948 , n21831 );
    not g9790 ( n15374 , n6140 );
    and g9791 ( n27107 , n17962 , n30059 );
    or g9792 ( n14263 , n31227 , n28744 );
    nor g9793 ( n22024 , n6681 , n27732 );
    xnor g9794 ( n25171 , n18708 , n11775 );
    or g9795 ( n18335 , n12316 , n12445 );
    not g9796 ( n26646 , n28590 );
    not g9797 ( n31524 , n6098 );
    or g9798 ( n18072 , n29451 , n16947 );
    xnor g9799 ( n21515 , n26317 , n9350 );
    and g9800 ( n28152 , n22661 , n19232 );
    xnor g9801 ( n31641 , n8931 , n15558 );
    not g9802 ( n15075 , n21521 );
    not g9803 ( n11863 , n10071 );
    and g9804 ( n31200 , n6247 , n18955 );
    or g9805 ( n6777 , n2243 , n8417 );
    or g9806 ( n20649 , n17227 , n7408 );
    or g9807 ( n14127 , n13580 , n20412 );
    xor g9808 ( n14241 , n15038 , n4185 );
    or g9809 ( n18539 , n965 , n30045 );
    or g9810 ( n29887 , n12918 , n28207 );
    xnor g9811 ( n24503 , n16109 , n30706 );
    or g9812 ( n31557 , n22133 , n279 );
    xnor g9813 ( n18515 , n3591 , n21603 );
    or g9814 ( n15375 , n19245 , n19928 );
    xnor g9815 ( n23387 , n21185 , n27805 );
    nor g9816 ( n24085 , n15793 , n28203 );
    or g9817 ( n9257 , n30000 , n18251 );
    nor g9818 ( n18326 , n17771 , n5273 );
    nor g9819 ( n10093 , n21629 , n20973 );
    not g9820 ( n28102 , n8947 );
    xnor g9821 ( n17402 , n18179 , n27847 );
    not g9822 ( n9286 , n28154 );
    or g9823 ( n210 , n7573 , n29149 );
    or g9824 ( n16062 , n24012 , n21378 );
    or g9825 ( n31844 , n12727 , n15253 );
    and g9826 ( n24060 , n3150 , n9811 );
    or g9827 ( n8272 , n14676 , n10100 );
    not g9828 ( n23484 , n3914 );
    xnor g9829 ( n1167 , n10597 , n9341 );
    not g9830 ( n30731 , n8808 );
    nor g9831 ( n31183 , n31204 , n8991 );
    xnor g9832 ( n8053 , n26006 , n27534 );
    nor g9833 ( n23077 , n5685 , n8670 );
    xnor g9834 ( n23165 , n2128 , n25734 );
    not g9835 ( n23294 , n22421 );
    nor g9836 ( n23334 , n12364 , n11416 );
    or g9837 ( n25275 , n27883 , n26002 );
    nor g9838 ( n14029 , n24776 , n15130 );
    and g9839 ( n22891 , n3704 , n20440 );
    xnor g9840 ( n13183 , n2695 , n17879 );
    not g9841 ( n29890 , n10978 );
    nor g9842 ( n540 , n1693 , n12603 );
    nor g9843 ( n16103 , n24794 , n31500 );
    xnor g9844 ( n14308 , n30831 , n11866 );
    xnor g9845 ( n2732 , n18901 , n14546 );
    or g9846 ( n27167 , n14325 , n29508 );
    xnor g9847 ( n20393 , n22519 , n4254 );
    or g9848 ( n11632 , n50 , n5013 );
    xnor g9849 ( n15835 , n16729 , n26496 );
    or g9850 ( n31064 , n1725 , n30994 );
    not g9851 ( n18688 , n16098 );
    xnor g9852 ( n24947 , n4765 , n24281 );
    and g9853 ( n15720 , n14068 , n26838 );
    or g9854 ( n18206 , n27877 , n19414 );
    or g9855 ( n2081 , n18263 , n7429 );
    and g9856 ( n18739 , n28906 , n4358 );
    not g9857 ( n11958 , n27355 );
    nor g9858 ( n15102 , n5136 , n4023 );
    nor g9859 ( n1647 , n31780 , n5990 );
    not g9860 ( n6760 , n21327 );
    not g9861 ( n26207 , n6140 );
    or g9862 ( n9919 , n8031 , n859 );
    and g9863 ( n1580 , n5802 , n19342 );
    and g9864 ( n23704 , n18937 , n9160 );
    xnor g9865 ( n454 , n11832 , n20295 );
    not g9866 ( n8966 , n11381 );
    not g9867 ( n26151 , n12849 );
    not g9868 ( n16835 , n7813 );
    xnor g9869 ( n6211 , n13699 , n14780 );
    or g9870 ( n31405 , n19001 , n7165 );
    and g9871 ( n9139 , n9104 , n26871 );
    or g9872 ( n22572 , n11789 , n28658 );
    xnor g9873 ( n20494 , n16859 , n26256 );
    xor g9874 ( n17808 , n7303 , n14847 );
    and g9875 ( n6690 , n6053 , n25778 );
    nor g9876 ( n25246 , n30287 , n2744 );
    not g9877 ( n22854 , n31474 );
    not g9878 ( n6070 , n21707 );
    or g9879 ( n9441 , n1450 , n16839 );
    or g9880 ( n27319 , n14157 , n7136 );
    not g9881 ( n25866 , n23595 );
    xnor g9882 ( n6754 , n6441 , n9949 );
    or g9883 ( n25713 , n24084 , n2166 );
    xnor g9884 ( n25057 , n26069 , n1388 );
    and g9885 ( n13512 , n208 , n4431 );
    xnor g9886 ( n19110 , n22557 , n431 );
    or g9887 ( n30995 , n31857 , n13212 );
    xnor g9888 ( n5443 , n11644 , n3784 );
    nor g9889 ( n13762 , n24650 , n24736 );
    not g9890 ( n15475 , n392 );
    xnor g9891 ( n13037 , n29142 , n30263 );
    or g9892 ( n4068 , n26187 , n29582 );
    and g9893 ( n6339 , n28138 , n15729 );
    not g9894 ( n10733 , n23038 );
    not g9895 ( n18168 , n12651 );
    xnor g9896 ( n27757 , n19513 , n1909 );
    and g9897 ( n12121 , n5657 , n23575 );
    or g9898 ( n14784 , n8675 , n26465 );
    not g9899 ( n3645 , n26657 );
    or g9900 ( n2229 , n7900 , n7172 );
    not g9901 ( n28411 , n16347 );
    xnor g9902 ( n29330 , n31141 , n1601 );
    not g9903 ( n23172 , n13868 );
    not g9904 ( n31865 , n22020 );
    and g9905 ( n8814 , n21483 , n5470 );
    not g9906 ( n19877 , n10507 );
    xnor g9907 ( n19106 , n17319 , n24601 );
    not g9908 ( n1453 , n10879 );
    or g9909 ( n22524 , n9069 , n11396 );
    or g9910 ( n2341 , n30405 , n29472 );
    xor g9911 ( n10759 , n16713 , n9509 );
    and g9912 ( n21927 , n16372 , n29058 );
    xnor g9913 ( n30337 , n13262 , n12794 );
    or g9914 ( n12560 , n27028 , n13499 );
    xnor g9915 ( n27648 , n4137 , n17048 );
    xnor g9916 ( n24734 , n12803 , n1057 );
    nor g9917 ( n3940 , n23023 , n26700 );
    not g9918 ( n31138 , n15064 );
    and g9919 ( n30570 , n19325 , n8001 );
    xnor g9920 ( n27736 , n24472 , n20730 );
    not g9921 ( n26396 , n3440 );
    and g9922 ( n9054 , n25854 , n22278 );
    xnor g9923 ( n21849 , n378 , n20676 );
    and g9924 ( n10061 , n8274 , n25758 );
    not g9925 ( n18778 , n154 );
    xnor g9926 ( n23689 , n21528 , n22954 );
    not g9927 ( n25999 , n11010 );
    not g9928 ( n14653 , n22177 );
    and g9929 ( n4205 , n9745 , n11488 );
    or g9930 ( n19135 , n15878 , n1508 );
    or g9931 ( n29128 , n30309 , n27810 );
    nor g9932 ( n29443 , n10490 , n12024 );
    xnor g9933 ( n14408 , n31111 , n26665 );
    or g9934 ( n22972 , n13736 , n21704 );
    xnor g9935 ( n16072 , n29542 , n17149 );
    xnor g9936 ( n23037 , n6075 , n13780 );
    not g9937 ( n7205 , n27034 );
    or g9938 ( n10777 , n22049 , n25247 );
    nor g9939 ( n11152 , n25332 , n5238 );
    or g9940 ( n14216 , n24712 , n8433 );
    not g9941 ( n19896 , n28185 );
    and g9942 ( n8035 , n15149 , n19589 );
    xnor g9943 ( n29182 , n1376 , n10858 );
    not g9944 ( n28143 , n13992 );
    or g9945 ( n971 , n26700 , n4361 );
    or g9946 ( n20259 , n23119 , n19999 );
    not g9947 ( n7951 , n23738 );
    nor g9948 ( n27404 , n29937 , n8482 );
    or g9949 ( n29523 , n6788 , n12995 );
    nor g9950 ( n10552 , n29444 , n15584 );
    xnor g9951 ( n9445 , n18868 , n3455 );
    not g9952 ( n32027 , n25228 );
    xnor g9953 ( n6114 , n29429 , n29454 );
    or g9954 ( n9409 , n21789 , n8576 );
    not g9955 ( n21369 , n1829 );
    or g9956 ( n16659 , n4038 , n16880 );
    xnor g9957 ( n29412 , n26901 , n29497 );
    not g9958 ( n24694 , n15365 );
    and g9959 ( n31097 , n30876 , n23084 );
    or g9960 ( n13428 , n19867 , n2817 );
    and g9961 ( n28195 , n3041 , n29278 );
    not g9962 ( n13629 , n7876 );
    not g9963 ( n7663 , n24132 );
    not g9964 ( n26997 , n25119 );
    and g9965 ( n15664 , n2128 , n25230 );
    not g9966 ( n24981 , n4262 );
    xnor g9967 ( n8874 , n11285 , n13404 );
    not g9968 ( n23177 , n22697 );
    and g9969 ( n4717 , n31893 , n9229 );
    nor g9970 ( n7654 , n24807 , n5339 );
    not g9971 ( n21961 , n16151 );
    not g9972 ( n4106 , n14838 );
    and g9973 ( n15861 , n14219 , n21210 );
    xnor g9974 ( n10902 , n23561 , n3268 );
    xnor g9975 ( n21356 , n12208 , n28727 );
    xnor g9976 ( n17781 , n11740 , n21708 );
    not g9977 ( n9029 , n21855 );
    or g9978 ( n8851 , n22843 , n2725 );
    and g9979 ( n10166 , n24688 , n19833 );
    xnor g9980 ( n1546 , n22184 , n3432 );
    xnor g9981 ( n8194 , n5625 , n9156 );
    not g9982 ( n12832 , n4107 );
    or g9983 ( n27277 , n12625 , n7619 );
    xor g9984 ( n3306 , n15279 , n27678 );
    or g9985 ( n30353 , n5603 , n2901 );
    not g9986 ( n3626 , n8185 );
    and g9987 ( n12083 , n12703 , n19592 );
    or g9988 ( n28743 , n27120 , n22815 );
    nor g9989 ( n28342 , n7596 , n22577 );
    and g9990 ( n20430 , n3705 , n25263 );
    not g9991 ( n14387 , n26087 );
    or g9992 ( n22957 , n26873 , n24601 );
    or g9993 ( n10384 , n9014 , n13863 );
    xnor g9994 ( n78 , n6619 , n29578 );
    not g9995 ( n16099 , n1484 );
    nor g9996 ( n13717 , n10548 , n20941 );
    xnor g9997 ( n20130 , n16659 , n21834 );
    or g9998 ( n19645 , n20524 , n16613 );
    not g9999 ( n14909 , n7709 );
    not g10000 ( n21010 , n27486 );
    not g10001 ( n27374 , n13514 );
    not g10002 ( n29401 , n8582 );
    not g10003 ( n7927 , n31543 );
    not g10004 ( n6428 , n17525 );
    not g10005 ( n31689 , n27690 );
    or g10006 ( n472 , n10474 , n5220 );
    xnor g10007 ( n17584 , n9921 , n7634 );
    or g10008 ( n26693 , n2290 , n3738 );
    not g10009 ( n28077 , n14807 );
    xnor g10010 ( n31857 , n25384 , n22177 );
    or g10011 ( n11083 , n8524 , n10406 );
    or g10012 ( n16588 , n4722 , n12677 );
    xnor g10013 ( n28854 , n19777 , n6370 );
    xnor g10014 ( n31323 , n28197 , n27625 );
    xor g10015 ( n9934 , n24495 , n9043 );
    buf g10016 ( n3182 , n18487 );
    xnor g10017 ( n13140 , n1313 , n10889 );
    or g10018 ( n17994 , n9011 , n2510 );
    or g10019 ( n10233 , n30133 , n27953 );
    not g10020 ( n18027 , n18889 );
    xnor g10021 ( n23692 , n25304 , n4367 );
    xnor g10022 ( n5187 , n19690 , n19379 );
    or g10023 ( n27592 , n8004 , n29252 );
    not g10024 ( n23948 , n22295 );
    xnor g10025 ( n12287 , n2820 , n22592 );
    xnor g10026 ( n10278 , n7820 , n494 );
    xor g10027 ( n20990 , n22127 , n20631 );
    not g10028 ( n25364 , n28212 );
    xnor g10029 ( n2906 , n445 , n26114 );
    and g10030 ( n5217 , n9245 , n22969 );
    not g10031 ( n22594 , n30801 );
    not g10032 ( n22710 , n24496 );
    not g10033 ( n11162 , n6801 );
    or g10034 ( n12854 , n25864 , n14507 );
    not g10035 ( n30658 , n10527 );
    not g10036 ( n21951 , n19939 );
    xor g10037 ( n9708 , n17547 , n2454 );
    or g10038 ( n10531 , n4732 , n18699 );
    not g10039 ( n9520 , n18391 );
    nor g10040 ( n25940 , n14035 , n3057 );
    not g10041 ( n26767 , n7722 );
    nor g10042 ( n14900 , n15987 , n27075 );
    and g10043 ( n24026 , n20460 , n5362 );
    or g10044 ( n31177 , n12806 , n25445 );
    or g10045 ( n28317 , n17229 , n1984 );
    nor g10046 ( n30902 , n29196 , n8114 );
    or g10047 ( n3127 , n25950 , n22044 );
    not g10048 ( n9147 , n9206 );
    not g10049 ( n12703 , n31868 );
    or g10050 ( n30914 , n25900 , n15557 );
    or g10051 ( n12907 , n19066 , n24712 );
    nor g10052 ( n21804 , n20825 , n1891 );
    xnor g10053 ( n9845 , n13376 , n19317 );
    xnor g10054 ( n16601 , n4816 , n13944 );
    or g10055 ( n29122 , n17368 , n31679 );
    and g10056 ( n17881 , n10816 , n18797 );
    or g10057 ( n15566 , n14424 , n1279 );
    or g10058 ( n29193 , n6145 , n26923 );
    and g10059 ( n14853 , n24403 , n25406 );
    not g10060 ( n9964 , n9669 );
    not g10061 ( n13471 , n25296 );
    and g10062 ( n26350 , n1060 , n30226 );
    nor g10063 ( n28810 , n19255 , n25115 );
    or g10064 ( n388 , n24917 , n26675 );
    not g10065 ( n25842 , n22379 );
    and g10066 ( n30946 , n4775 , n17999 );
    not g10067 ( n19702 , n4316 );
    xnor g10068 ( n5957 , n18791 , n391 );
    not g10069 ( n11288 , n28617 );
    not g10070 ( n1354 , n15425 );
    nor g10071 ( n7793 , n13579 , n470 );
    nor g10072 ( n1305 , n21261 , n14413 );
    or g10073 ( n22092 , n24830 , n2134 );
    not g10074 ( n30852 , n27210 );
    or g10075 ( n24529 , n28174 , n29602 );
    or g10076 ( n31298 , n18051 , n28429 );
    or g10077 ( n29943 , n31722 , n16711 );
    not g10078 ( n18462 , n142 );
    or g10079 ( n635 , n20608 , n1006 );
    and g10080 ( n5745 , n14797 , n21734 );
    or g10081 ( n30760 , n23354 , n14103 );
    or g10082 ( n27699 , n8597 , n3516 );
    xnor g10083 ( n14175 , n29569 , n24066 );
    xnor g10084 ( n8449 , n18353 , n20653 );
    nor g10085 ( n30949 , n6935 , n14514 );
    xnor g10086 ( n29620 , n16558 , n7046 );
    xnor g10087 ( n27432 , n9240 , n16594 );
    xor g10088 ( n5003 , n16087 , n23902 );
    xnor g10089 ( n981 , n14468 , n10370 );
    nor g10090 ( n26718 , n8988 , n30676 );
    and g10091 ( n5061 , n12675 , n16454 );
    and g10092 ( n15116 , n27399 , n29512 );
    not g10093 ( n27420 , n26269 );
    or g10094 ( n27843 , n23811 , n2689 );
    nor g10095 ( n13418 , n11645 , n30418 );
    or g10096 ( n23072 , n21371 , n15975 );
    xnor g10097 ( n11840 , n20609 , n8977 );
    xnor g10098 ( n30513 , n7939 , n12024 );
    not g10099 ( n24 , n18339 );
    or g10100 ( n6157 , n20532 , n19760 );
    and g10101 ( n15249 , n8834 , n23040 );
    and g10102 ( n8258 , n14156 , n28485 );
    or g10103 ( n429 , n3036 , n15620 );
    nor g10104 ( n12691 , n17068 , n18157 );
    nor g10105 ( n23114 , n10532 , n6905 );
    or g10106 ( n21046 , n30002 , n9655 );
    or g10107 ( n29175 , n12035 , n4359 );
    or g10108 ( n1926 , n20846 , n12477 );
    and g10109 ( n31068 , n26214 , n13597 );
    or g10110 ( n11186 , n20664 , n1632 );
    or g10111 ( n380 , n20417 , n12100 );
    xnor g10112 ( n16008 , n25845 , n5641 );
    and g10113 ( n16344 , n30930 , n16483 );
    xnor g10114 ( n24456 , n28950 , n19114 );
    not g10115 ( n28521 , n13886 );
    or g10116 ( n20592 , n35 , n11242 );
    not g10117 ( n596 , n7209 );
    buf g10118 ( n11257 , n17713 );
    xnor g10119 ( n14996 , n28913 , n8919 );
    not g10120 ( n4022 , n21015 );
    and g10121 ( n4340 , n3739 , n6037 );
    xnor g10122 ( n8400 , n26399 , n9873 );
    or g10123 ( n16243 , n14010 , n18023 );
    not g10124 ( n21851 , n26047 );
    or g10125 ( n9823 , n4640 , n13967 );
    xnor g10126 ( n13012 , n18465 , n23708 );
    or g10127 ( n26143 , n17706 , n15953 );
    xnor g10128 ( n17952 , n20010 , n17054 );
    not g10129 ( n653 , n14690 );
    xnor g10130 ( n18691 , n15131 , n18382 );
    xnor g10131 ( n13402 , n26074 , n29289 );
    or g10132 ( n25863 , n28433 , n22383 );
    xnor g10133 ( n22207 , n20550 , n30656 );
    not g10134 ( n18606 , n25415 );
    not g10135 ( n4002 , n25757 );
    not g10136 ( n25093 , n29587 );
    or g10137 ( n30834 , n20902 , n12938 );
    nor g10138 ( n8794 , n17517 , n29157 );
    and g10139 ( n19822 , n24264 , n6417 );
    xnor g10140 ( n1008 , n5891 , n7942 );
    not g10141 ( n4922 , n28741 );
    not g10142 ( n6355 , n19083 );
    not g10143 ( n11668 , n14214 );
    and g10144 ( n14327 , n10993 , n9102 );
    and g10145 ( n3260 , n22791 , n7015 );
    or g10146 ( n23465 , n10138 , n19123 );
    not g10147 ( n12355 , n25701 );
    and g10148 ( n21821 , n24619 , n11544 );
    or g10149 ( n6854 , n25276 , n4629 );
    or g10150 ( n29325 , n21603 , n30553 );
    or g10151 ( n1739 , n20365 , n24335 );
    not g10152 ( n4923 , n1755 );
    xnor g10153 ( n13615 , n658 , n17474 );
    not g10154 ( n14735 , n27769 );
    or g10155 ( n16143 , n1839 , n15684 );
    or g10156 ( n5070 , n19537 , n6095 );
    xnor g10157 ( n13237 , n31841 , n14316 );
    xnor g10158 ( n20170 , n19402 , n2851 );
    not g10159 ( n31561 , n2235 );
    and g10160 ( n30080 , n30234 , n30112 );
    not g10161 ( n17162 , n15132 );
    not g10162 ( n23556 , n24305 );
    or g10163 ( n1937 , n16921 , n26742 );
    not g10164 ( n19399 , n14451 );
    not g10165 ( n30754 , n15829 );
    not g10166 ( n18753 , n17441 );
    xnor g10167 ( n1786 , n1942 , n4393 );
    or g10168 ( n11773 , n10074 , n14590 );
    xnor g10169 ( n13812 , n30629 , n346 );
    nor g10170 ( n3158 , n10135 , n9556 );
    not g10171 ( n16732 , n23626 );
    not g10172 ( n23533 , n28674 );
    or g10173 ( n9620 , n13988 , n13541 );
    not g10174 ( n24355 , n13501 );
    or g10175 ( n13931 , n554 , n7514 );
    or g10176 ( n27007 , n21693 , n23923 );
    xnor g10177 ( n18676 , n31431 , n5975 );
    or g10178 ( n27603 , n21910 , n21955 );
    or g10179 ( n1747 , n9604 , n21521 );
    xnor g10180 ( n31981 , n24768 , n5723 );
    xnor g10181 ( n20891 , n2077 , n11937 );
    and g10182 ( n20829 , n25853 , n7631 );
    or g10183 ( n24755 , n16489 , n20399 );
    not g10184 ( n9518 , n6818 );
    nor g10185 ( n25147 , n10922 , n21249 );
    not g10186 ( n24110 , n11392 );
    not g10187 ( n8995 , n7583 );
    xnor g10188 ( n27681 , n14477 , n21136 );
    buf g10189 ( n22870 , n24703 );
    or g10190 ( n9364 , n20970 , n15972 );
    xnor g10191 ( n2986 , n11852 , n28828 );
    not g10192 ( n8290 , n27454 );
    xnor g10193 ( n24089 , n20309 , n20050 );
    not g10194 ( n29413 , n19826 );
    and g10195 ( n24856 , n1047 , n23933 );
    and g10196 ( n18088 , n22343 , n10914 );
    or g10197 ( n25921 , n27073 , n31242 );
    xnor g10198 ( n15822 , n15080 , n20575 );
    or g10199 ( n31059 , n19257 , n20090 );
    xnor g10200 ( n12942 , n27167 , n14469 );
    xnor g10201 ( n22218 , n4734 , n21890 );
    nor g10202 ( n12676 , n22349 , n25405 );
    not g10203 ( n5772 , n30856 );
    and g10204 ( n6234 , n23849 , n30952 );
    not g10205 ( n15936 , n10883 );
    xnor g10206 ( n26678 , n22841 , n9744 );
    not g10207 ( n20548 , n1145 );
    xnor g10208 ( n16334 , n22365 , n22016 );
    xnor g10209 ( n12255 , n22545 , n2559 );
    and g10210 ( n9677 , n4655 , n20354 );
    not g10211 ( n9940 , n31634 );
    not g10212 ( n20573 , n18017 );
    or g10213 ( n6638 , n6486 , n161 );
    xnor g10214 ( n12911 , n15299 , n6556 );
    or g10215 ( n29256 , n16759 , n2799 );
    not g10216 ( n1615 , n1877 );
    nor g10217 ( n7183 , n14732 , n10908 );
    xnor g10218 ( n16288 , n30302 , n19316 );
    and g10219 ( n26766 , n1851 , n17858 );
    not g10220 ( n8838 , n22169 );
    or g10221 ( n17359 , n27276 , n12091 );
    or g10222 ( n29046 , n1182 , n16556 );
    xnor g10223 ( n228 , n3892 , n2578 );
    xnor g10224 ( n1676 , n25173 , n20111 );
    xnor g10225 ( n21781 , n2917 , n25177 );
    or g10226 ( n4639 , n86 , n18158 );
    and g10227 ( n30550 , n27874 , n24186 );
    nor g10228 ( n30561 , n21485 , n23232 );
    and g10229 ( n2423 , n29328 , n5976 );
    and g10230 ( n30841 , n25951 , n7069 );
    nor g10231 ( n16892 , n6641 , n22943 );
    and g10232 ( n5433 , n31967 , n17850 );
    not g10233 ( n27486 , n12788 );
    not g10234 ( n1035 , n18907 );
    and g10235 ( n52 , n22072 , n25024 );
    or g10236 ( n28669 , n11990 , n5304 );
    or g10237 ( n28038 , n31896 , n12479 );
    or g10238 ( n21451 , n1358 , n5455 );
    not g10239 ( n19768 , n6739 );
    buf g10240 ( n5559 , n28209 );
    or g10241 ( n31219 , n1148 , n4440 );
    xnor g10242 ( n18246 , n16222 , n30525 );
    not g10243 ( n30459 , n3568 );
    not g10244 ( n7855 , n20400 );
    xnor g10245 ( n13974 , n20054 , n15464 );
    not g10246 ( n7157 , n13124 );
    xnor g10247 ( n23802 , n4184 , n17781 );
    buf g10248 ( n27995 , n3276 );
    not g10249 ( n31310 , n9190 );
    not g10250 ( n26308 , n27215 );
    and g10251 ( n10596 , n13240 , n22348 );
    xnor g10252 ( n30084 , n24118 , n28983 );
    xnor g10253 ( n29109 , n28397 , n14136 );
    xnor g10254 ( n1 , n10164 , n27949 );
    and g10255 ( n20302 , n31833 , n1459 );
    xnor g10256 ( n21008 , n26654 , n16308 );
    xnor g10257 ( n16403 , n22637 , n28445 );
    and g10258 ( n1833 , n29842 , n346 );
    nor g10259 ( n13669 , n7314 , n6191 );
    xnor g10260 ( n29932 , n8121 , n5297 );
    not g10261 ( n31835 , n20120 );
    xnor g10262 ( n4943 , n24158 , n8931 );
    and g10263 ( n25360 , n7347 , n29866 );
    and g10264 ( n30215 , n5103 , n8567 );
    or g10265 ( n12565 , n4554 , n228 );
    or g10266 ( n1079 , n11473 , n16354 );
    or g10267 ( n9593 , n17877 , n25426 );
    not g10268 ( n30145 , n17928 );
    xnor g10269 ( n29129 , n13093 , n10917 );
    not g10270 ( n14359 , n18889 );
    xnor g10271 ( n3382 , n9114 , n19855 );
    and g10272 ( n27941 , n46 , n27968 );
    not g10273 ( n17954 , n4375 );
    xnor g10274 ( n5523 , n19230 , n11778 );
    not g10275 ( n18669 , n1545 );
    or g10276 ( n9630 , n29105 , n8027 );
    xor g10277 ( n29435 , n22789 , n24761 );
    and g10278 ( n25228 , n28775 , n5283 );
    not g10279 ( n21244 , n3845 );
    xnor g10280 ( n8158 , n29217 , n22045 );
    xnor g10281 ( n18672 , n8899 , n13293 );
    and g10282 ( n23641 , n20690 , n12933 );
    or g10283 ( n22771 , n14398 , n21509 );
    or g10284 ( n18013 , n107 , n20600 );
    xnor g10285 ( n23378 , n25183 , n24466 );
    not g10286 ( n394 , n16722 );
    and g10287 ( n9550 , n30032 , n22356 );
    and g10288 ( n12661 , n24489 , n28013 );
    and g10289 ( n7774 , n7169 , n31047 );
    not g10290 ( n9856 , n1322 );
    or g10291 ( n10567 , n15897 , n18644 );
    or g10292 ( n11403 , n26114 , n30046 );
    xnor g10293 ( n13380 , n19618 , n324 );
    and g10294 ( n15209 , n25191 , n27277 );
    or g10295 ( n22969 , n30074 , n6739 );
    and g10296 ( n25477 , n1094 , n12147 );
    or g10297 ( n23146 , n8707 , n26578 );
    xnor g10298 ( n21733 , n12914 , n21028 );
    xnor g10299 ( n14456 , n22731 , n16381 );
    nor g10300 ( n13825 , n16300 , n27615 );
    not g10301 ( n29217 , n20842 );
    and g10302 ( n29026 , n22132 , n14294 );
    not g10303 ( n23391 , n11424 );
    and g10304 ( n17315 , n29009 , n15046 );
    xnor g10305 ( n13959 , n5388 , n9509 );
    xnor g10306 ( n18090 , n23921 , n30498 );
    or g10307 ( n14587 , n7315 , n28632 );
    not g10308 ( n15586 , n11220 );
    xnor g10309 ( n29073 , n1239 , n17207 );
    nor g10310 ( n10409 , n16132 , n25668 );
    and g10311 ( n9038 , n11448 , n30206 );
    or g10312 ( n5920 , n1775 , n27826 );
    xnor g10313 ( n21402 , n674 , n320 );
    not g10314 ( n11247 , n1670 );
    and g10315 ( n23805 , n8828 , n13929 );
    or g10316 ( n25464 , n31727 , n30585 );
    xnor g10317 ( n32004 , n3885 , n21679 );
    nor g10318 ( n22010 , n3631 , n19991 );
    not g10319 ( n31819 , n19333 );
    or g10320 ( n17314 , n13008 , n30965 );
    or g10321 ( n18020 , n28283 , n26954 );
    and g10322 ( n8954 , n22337 , n13009 );
    not g10323 ( n19754 , n7180 );
    not g10324 ( n1194 , n4149 );
    and g10325 ( n6275 , n5034 , n15922 );
    xnor g10326 ( n22592 , n28033 , n27742 );
    not g10327 ( n12812 , n26279 );
    and g10328 ( n3245 , n6937 , n11281 );
    and g10329 ( n31004 , n5104 , n20867 );
    or g10330 ( n31612 , n5222 , n25280 );
    or g10331 ( n23028 , n6999 , n3374 );
    not g10332 ( n21425 , n2022 );
    not g10333 ( n13155 , n25007 );
    not g10334 ( n24765 , n3276 );
    not g10335 ( n26555 , n14040 );
    xnor g10336 ( n27789 , n13024 , n2673 );
    or g10337 ( n19863 , n6690 , n11503 );
    or g10338 ( n9452 , n28748 , n6245 );
    xnor g10339 ( n23365 , n12724 , n19632 );
    or g10340 ( n11418 , n4045 , n20864 );
    not g10341 ( n22174 , n1010 );
    not g10342 ( n29629 , n4397 );
    or g10343 ( n3272 , n20865 , n24008 );
    and g10344 ( n26160 , n28456 , n2419 );
    not g10345 ( n11796 , n9334 );
    xnor g10346 ( n4218 , n24074 , n10921 );
    not g10347 ( n28258 , n21597 );
    xnor g10348 ( n17914 , n29726 , n26615 );
    not g10349 ( n19404 , n1999 );
    not g10350 ( n20211 , n24487 );
    and g10351 ( n20752 , n25863 , n8123 );
    or g10352 ( n30475 , n29331 , n6032 );
    nor g10353 ( n7170 , n17254 , n9973 );
    and g10354 ( n22467 , n20981 , n3289 );
    xnor g10355 ( n5643 , n14349 , n12745 );
    or g10356 ( n24684 , n21731 , n2943 );
    not g10357 ( n24433 , n3804 );
    and g10358 ( n8127 , n2013 , n30066 );
    or g10359 ( n27563 , n26804 , n6335 );
    xnor g10360 ( n1241 , n6587 , n18908 );
    and g10361 ( n16615 , n23818 , n6184 );
    nor g10362 ( n8219 , n22755 , n26995 );
    or g10363 ( n14347 , n6583 , n10767 );
    or g10364 ( n18987 , n18342 , n30302 );
    not g10365 ( n18197 , n29601 );
    not g10366 ( n13779 , n12210 );
    not g10367 ( n22431 , n27092 );
    xnor g10368 ( n13219 , n11922 , n29490 );
    not g10369 ( n18311 , n19920 );
    xnor g10370 ( n22826 , n22610 , n25766 );
    or g10371 ( n25803 , n27343 , n24362 );
    nor g10372 ( n21681 , n2798 , n6374 );
    not g10373 ( n20877 , n13555 );
    and g10374 ( n17223 , n31642 , n15565 );
    or g10375 ( n18782 , n23572 , n11729 );
    xnor g10376 ( n19400 , n9347 , n4953 );
    or g10377 ( n12824 , n24066 , n4994 );
    or g10378 ( n8615 , n7803 , n6941 );
    not g10379 ( n11903 , n17924 );
    and g10380 ( n26059 , n29299 , n10424 );
    and g10381 ( n6062 , n1492 , n13490 );
    and g10382 ( n6506 , n5516 , n15032 );
    or g10383 ( n2594 , n30348 , n22438 );
    xnor g10384 ( n18025 , n11732 , n25513 );
    xnor g10385 ( n5862 , n20971 , n9424 );
    xnor g10386 ( n4107 , n7173 , n24004 );
    or g10387 ( n4236 , n5783 , n31435 );
    not g10388 ( n4277 , n9339 );
    nor g10389 ( n15896 , n11197 , n30412 );
    xnor g10390 ( n18012 , n28651 , n31020 );
    and g10391 ( n4858 , n26935 , n19544 );
    or g10392 ( n15032 , n13421 , n18337 );
    or g10393 ( n1874 , n25866 , n28718 );
    not g10394 ( n2244 , n21165 );
    and g10395 ( n13988 , n11434 , n15192 );
    and g10396 ( n26634 , n27378 , n15353 );
    and g10397 ( n19815 , n7271 , n27838 );
    and g10398 ( n3135 , n12471 , n9604 );
    xnor g10399 ( n24037 , n16531 , n17125 );
    and g10400 ( n2514 , n28658 , n11789 );
    nor g10401 ( n7158 , n9011 , n14112 );
    and g10402 ( n19758 , n7523 , n23592 );
    not g10403 ( n4428 , n891 );
    not g10404 ( n3203 , n25042 );
    not g10405 ( n14770 , n9524 );
    and g10406 ( n10382 , n954 , n7601 );
    not g10407 ( n11859 , n24268 );
    not g10408 ( n3284 , n29829 );
    not g10409 ( n24546 , n4686 );
    or g10410 ( n11114 , n25806 , n16698 );
    not g10411 ( n3004 , n14290 );
    xnor g10412 ( n31278 , n2540 , n18259 );
    xnor g10413 ( n26683 , n23155 , n8222 );
    not g10414 ( n10748 , n5768 );
    xnor g10415 ( n24163 , n16569 , n22075 );
    not g10416 ( n15357 , n24914 );
    nor g10417 ( n9808 , n10477 , n13918 );
    not g10418 ( n10589 , n13329 );
    not g10419 ( n10291 , n1166 );
    xnor g10420 ( n14003 , n7679 , n17304 );
    and g10421 ( n6600 , n7716 , n16917 );
    or g10422 ( n2534 , n15824 , n27861 );
    not g10423 ( n14882 , n8853 );
    xnor g10424 ( n26094 , n27953 , n10736 );
    and g10425 ( n23594 , n21325 , n27284 );
    not g10426 ( n9627 , n4560 );
    not g10427 ( n7919 , n1099 );
    not g10428 ( n19652 , n18831 );
    or g10429 ( n6033 , n7565 , n17741 );
    not g10430 ( n12639 , n13649 );
    xnor g10431 ( n14837 , n9438 , n22796 );
    nor g10432 ( n4545 , n15999 , n1100 );
    not g10433 ( n21581 , n19959 );
    xnor g10434 ( n30285 , n20759 , n28634 );
    xnor g10435 ( n19359 , n29390 , n14954 );
    not g10436 ( n14093 , n26795 );
    or g10437 ( n23425 , n1089 , n19290 );
    or g10438 ( n32015 , n30044 , n27652 );
    xor g10439 ( n20531 , n27992 , n14473 );
    not g10440 ( n8893 , n10032 );
    xnor g10441 ( n22412 , n470 , n1692 );
    buf g10442 ( n16299 , n18322 );
    not g10443 ( n8947 , n11286 );
    xnor g10444 ( n6412 , n31752 , n15266 );
    and g10445 ( n31149 , n18579 , n27387 );
    xnor g10446 ( n5986 , n24249 , n12546 );
    xnor g10447 ( n29372 , n19702 , n11281 );
    xnor g10448 ( n12135 , n4364 , n27849 );
    and g10449 ( n21922 , n15765 , n6501 );
    and g10450 ( n6767 , n8049 , n5858 );
    nor g10451 ( n27793 , n15178 , n21926 );
    or g10452 ( n30665 , n8561 , n13343 );
    not g10453 ( n23417 , n25436 );
    or g10454 ( n26721 , n12312 , n10346 );
    nor g10455 ( n12144 , n17310 , n21225 );
    or g10456 ( n30499 , n5704 , n30959 );
    or g10457 ( n14804 , n21233 , n7650 );
    not g10458 ( n6751 , n31002 );
    xnor g10459 ( n29045 , n10446 , n12082 );
    and g10460 ( n26493 , n30901 , n25597 );
    xnor g10461 ( n25438 , n14555 , n31019 );
    not g10462 ( n26212 , n16654 );
    and g10463 ( n31096 , n14784 , n10915 );
    not g10464 ( n18900 , n12817 );
    or g10465 ( n28813 , n26598 , n3698 );
    or g10466 ( n27423 , n29667 , n7651 );
    xnor g10467 ( n6801 , n15396 , n614 );
    not g10468 ( n5868 , n11425 );
    or g10469 ( n2772 , n7014 , n12170 );
    xnor g10470 ( n8689 , n30123 , n5555 );
    xnor g10471 ( n7962 , n13254 , n22251 );
    nor g10472 ( n23240 , n6495 , n30806 );
    and g10473 ( n25985 , n17708 , n23822 );
    xnor g10474 ( n29838 , n17897 , n13299 );
    xnor g10475 ( n20407 , n17605 , n30338 );
    not g10476 ( n16033 , n21300 );
    nor g10477 ( n28682 , n6166 , n9300 );
    or g10478 ( n23272 , n27536 , n27089 );
    buf g10479 ( n27546 , n20251 );
    or g10480 ( n11165 , n18413 , n190 );
    xnor g10481 ( n14484 , n18971 , n31540 );
    or g10482 ( n30299 , n28392 , n21739 );
    xnor g10483 ( n30670 , n14670 , n7465 );
    or g10484 ( n22889 , n23476 , n6515 );
    xnor g10485 ( n6525 , n8497 , n12777 );
    and g10486 ( n27246 , n25969 , n1874 );
    xnor g10487 ( n23885 , n10379 , n15838 );
    not g10488 ( n2068 , n6524 );
    not g10489 ( n5836 , n25366 );
    xnor g10490 ( n16522 , n29971 , n22456 );
    and g10491 ( n16931 , n13033 , n20301 );
    and g10492 ( n16727 , n6795 , n30726 );
    and g10493 ( n28450 , n26787 , n31773 );
    nor g10494 ( n12095 , n21464 , n13319 );
    xnor g10495 ( n1010 , n24091 , n22475 );
    or g10496 ( n18927 , n15337 , n5325 );
    xnor g10497 ( n27658 , n24170 , n28514 );
    xnor g10498 ( n31505 , n26646 , n16762 );
    or g10499 ( n3129 , n27708 , n17616 );
    or g10500 ( n9687 , n13801 , n30216 );
    nor g10501 ( n15173 , n26894 , n6874 );
    nor g10502 ( n30344 , n30467 , n10194 );
    or g10503 ( n12823 , n7584 , n17345 );
    xnor g10504 ( n13826 , n1643 , n11617 );
    xnor g10505 ( n15293 , n23230 , n11110 );
    not g10506 ( n25591 , n19250 );
    not g10507 ( n218 , n23045 );
    not g10508 ( n22124 , n17790 );
    nor g10509 ( n5130 , n12668 , n13680 );
    not g10510 ( n31034 , n29010 );
    xnor g10511 ( n22757 , n29842 , n346 );
    xnor g10512 ( n9703 , n7748 , n17194 );
    xor g10513 ( n17509 , n5806 , n2288 );
    nor g10514 ( n11479 , n10119 , n10716 );
    and g10515 ( n14281 , n9704 , n28842 );
    or g10516 ( n28454 , n13727 , n8974 );
    not g10517 ( n25972 , n20692 );
    or g10518 ( n2020 , n26627 , n15044 );
    xnor g10519 ( n20976 , n10777 , n19793 );
    or g10520 ( n9841 , n23162 , n22288 );
    and g10521 ( n30397 , n9995 , n28493 );
    or g10522 ( n24906 , n823 , n1994 );
    or g10523 ( n24801 , n4046 , n9191 );
    xnor g10524 ( n11719 , n23040 , n17255 );
    nor g10525 ( n21888 , n4257 , n11262 );
    xnor g10526 ( n31073 , n9243 , n6830 );
    not g10527 ( n10934 , n14336 );
    xnor g10528 ( n553 , n6691 , n31888 );
    xnor g10529 ( n18512 , n12270 , n20129 );
    not g10530 ( n18189 , n7894 );
    nor g10531 ( n4084 , n2862 , n3432 );
    not g10532 ( n10125 , n18857 );
    xnor g10533 ( n7455 , n7718 , n28081 );
    or g10534 ( n10575 , n20944 , n2011 );
    nor g10535 ( n9281 , n14488 , n6278 );
    xnor g10536 ( n2204 , n19736 , n6489 );
    or g10537 ( n273 , n24584 , n23776 );
    or g10538 ( n29465 , n21687 , n28151 );
    not g10539 ( n2938 , n28384 );
    nor g10540 ( n25113 , n18389 , n4213 );
    or g10541 ( n17373 , n12492 , n576 );
    not g10542 ( n23179 , n3907 );
    xnor g10543 ( n5362 , n283 , n13437 );
    not g10544 ( n6697 , n31928 );
    xnor g10545 ( n6184 , n16420 , n20865 );
    or g10546 ( n11027 , n27807 , n22056 );
    xor g10547 ( n26284 , n21406 , n29021 );
    not g10548 ( n13243 , n10981 );
    xnor g10549 ( n15074 , n26157 , n16055 );
    not g10550 ( n9349 , n13417 );
    or g10551 ( n13051 , n1670 , n16045 );
    not g10552 ( n30501 , n4624 );
    not g10553 ( n20186 , n17941 );
    xnor g10554 ( n30470 , n3822 , n23097 );
    nor g10555 ( n6716 , n1177 , n31470 );
    and g10556 ( n8748 , n27109 , n21272 );
    or g10557 ( n6197 , n7894 , n22650 );
    and g10558 ( n23772 , n28893 , n20838 );
    nor g10559 ( n23229 , n29902 , n10534 );
    xnor g10560 ( n21908 , n29939 , n18333 );
    and g10561 ( n15690 , n29564 , n14481 );
    or g10562 ( n18129 , n19472 , n8056 );
    not g10563 ( n4944 , n12759 );
    not g10564 ( n2728 , n30603 );
    not g10565 ( n9778 , n19340 );
    and g10566 ( n22630 , n1668 , n27891 );
    xnor g10567 ( n627 , n20434 , n9601 );
    not g10568 ( n7594 , n9766 );
    not g10569 ( n23673 , n6406 );
    or g10570 ( n16469 , n18086 , n444 );
    xnor g10571 ( n20801 , n349 , n13037 );
    xnor g10572 ( n14830 , n5865 , n24217 );
    and g10573 ( n29909 , n21097 , n1697 );
    and g10574 ( n23920 , n8121 , n23107 );
    and g10575 ( n6175 , n7842 , n4975 );
    not g10576 ( n29929 , n11947 );
    not g10577 ( n24644 , n3938 );
    or g10578 ( n7817 , n11934 , n28498 );
    or g10579 ( n8955 , n28828 , n19810 );
    nor g10580 ( n27654 , n26974 , n10676 );
    and g10581 ( n25279 , n19951 , n13191 );
    and g10582 ( n5861 , n20627 , n2290 );
    not g10583 ( n21610 , n4439 );
    xnor g10584 ( n2210 , n4865 , n16536 );
    and g10585 ( n104 , n11914 , n24928 );
    or g10586 ( n24597 , n3295 , n5814 );
    and g10587 ( n3130 , n8499 , n11297 );
    and g10588 ( n8930 , n6292 , n8243 );
    xnor g10589 ( n5728 , n5474 , n16998 );
    not g10590 ( n4096 , n27963 );
    not g10591 ( n2477 , n3443 );
    not g10592 ( n1375 , n22451 );
    xnor g10593 ( n10522 , n24304 , n29059 );
    and g10594 ( n10595 , n24953 , n31940 );
    or g10595 ( n20609 , n24257 , n22739 );
    not g10596 ( n4602 , n13708 );
    not g10597 ( n8207 , n3430 );
    and g10598 ( n18397 , n24821 , n13465 );
    or g10599 ( n24103 , n21308 , n23710 );
    xnor g10600 ( n6138 , n20664 , n31470 );
    not g10601 ( n2270 , n26510 );
    and g10602 ( n26102 , n10347 , n26523 );
    xnor g10603 ( n29369 , n15898 , n28166 );
    or g10604 ( n21397 , n11301 , n29431 );
    not g10605 ( n22523 , n31358 );
    xnor g10606 ( n8900 , n23597 , n16986 );
    xor g10607 ( n4000 , n24523 , n17649 );
    not g10608 ( n7716 , n24724 );
    and g10609 ( n17216 , n9233 , n30935 );
    not g10610 ( n31801 , n996 );
    and g10611 ( n30053 , n22303 , n18013 );
    not g10612 ( n31843 , n27487 );
    and g10613 ( n25281 , n4731 , n29174 );
    and g10614 ( n7245 , n6932 , n8992 );
    or g10615 ( n3434 , n6072 , n14100 );
    xnor g10616 ( n13591 , n21505 , n28958 );
    xnor g10617 ( n4266 , n24728 , n1236 );
    not g10618 ( n27955 , n8057 );
    xnor g10619 ( n18101 , n6227 , n30329 );
    or g10620 ( n22764 , n2447 , n6141 );
    xor g10621 ( n5338 , n11580 , n22845 );
    or g10622 ( n25514 , n28267 , n6651 );
    or g10623 ( n29480 , n29897 , n23321 );
    nor g10624 ( n7997 , n11785 , n975 );
    xnor g10625 ( n16653 , n13070 , n11702 );
    xnor g10626 ( n5697 , n24075 , n25123 );
    or g10627 ( n2084 , n30731 , n12978 );
    xnor g10628 ( n3783 , n2665 , n19632 );
    not g10629 ( n21233 , n4252 );
    and g10630 ( n16746 , n4365 , n3574 );
    and g10631 ( n27300 , n29233 , n23675 );
    or g10632 ( n29598 , n10383 , n7928 );
    or g10633 ( n2421 , n9915 , n1697 );
    xnor g10634 ( n1345 , n19683 , n24276 );
    nor g10635 ( n11274 , n365 , n13952 );
    not g10636 ( n13714 , n3315 );
    nor g10637 ( n16383 , n24525 , n1414 );
    xnor g10638 ( n25213 , n1054 , n7690 );
    not g10639 ( n17145 , n10091 );
    or g10640 ( n16590 , n3167 , n17252 );
    not g10641 ( n14567 , n6213 );
    xnor g10642 ( n13577 , n1061 , n3199 );
    not g10643 ( n2078 , n5685 );
    not g10644 ( n20484 , n17722 );
    not g10645 ( n19786 , n27443 );
    xnor g10646 ( n28075 , n3749 , n2861 );
    not g10647 ( n4807 , n1109 );
    not g10648 ( n3984 , n22550 );
    or g10649 ( n28118 , n30002 , n14566 );
    or g10650 ( n8165 , n26088 , n8258 );
    and g10651 ( n18478 , n4787 , n24375 );
    and g10652 ( n19703 , n13099 , n5366 );
    and g10653 ( n25076 , n7577 , n23496 );
    not g10654 ( n5909 , n171 );
    xnor g10655 ( n8718 , n29600 , n28806 );
    or g10656 ( n16235 , n12142 , n11774 );
    and g10657 ( n28723 , n15339 , n22772 );
    xnor g10658 ( n1335 , n29974 , n12035 );
    or g10659 ( n24922 , n29477 , n4460 );
    xnor g10660 ( n12617 , n8578 , n1983 );
    or g10661 ( n18276 , n24962 , n1799 );
    or g10662 ( n26304 , n2685 , n22168 );
    or g10663 ( n22330 , n16033 , n21113 );
    or g10664 ( n10132 , n18765 , n27729 );
    xnor g10665 ( n29862 , n31275 , n19212 );
    not g10666 ( n14960 , n5706 );
    nor g10667 ( n14264 , n26315 , n13743 );
    xnor g10668 ( n26302 , n18303 , n16468 );
    or g10669 ( n20197 , n1720 , n28440 );
    xnor g10670 ( n22348 , n5775 , n31428 );
    not g10671 ( n29036 , n9862 );
    or g10672 ( n24507 , n14329 , n29995 );
    or g10673 ( n25075 , n10671 , n14327 );
    nor g10674 ( n14767 , n26456 , n8042 );
    not g10675 ( n19025 , n31176 );
    not g10676 ( n3975 , n1995 );
    or g10677 ( n18075 , n332 , n29594 );
    and g10678 ( n25226 , n12370 , n20175 );
    and g10679 ( n27799 , n11427 , n27668 );
    not g10680 ( n6820 , n9948 );
    and g10681 ( n28573 , n3891 , n12869 );
    not g10682 ( n11458 , n16444 );
    xnor g10683 ( n5168 , n30297 , n10327 );
    and g10684 ( n25017 , n6321 , n29179 );
    not g10685 ( n7318 , n7562 );
    not g10686 ( n2644 , n6036 );
    not g10687 ( n21940 , n30281 );
    or g10688 ( n19116 , n25707 , n9911 );
    xnor g10689 ( n27403 , n22508 , n29421 );
    and g10690 ( n1150 , n31992 , n22350 );
    xnor g10691 ( n5588 , n19023 , n8399 );
    and g10692 ( n2035 , n665 , n18591 );
    and g10693 ( n24376 , n8659 , n27990 );
    xnor g10694 ( n784 , n26029 , n18955 );
    not g10695 ( n24040 , n1755 );
    not g10696 ( n14237 , n26364 );
    xnor g10697 ( n16080 , n8420 , n5122 );
    not g10698 ( n13791 , n11810 );
    not g10699 ( n9434 , n13397 );
    xnor g10700 ( n26422 , n6278 , n15010 );
    and g10701 ( n25116 , n7332 , n26071 );
    nor g10702 ( n11749 , n19078 , n26265 );
    buf g10703 ( n20278 , n31915 );
    and g10704 ( n27535 , n11590 , n8901 );
    or g10705 ( n7153 , n16132 , n5833 );
    xnor g10706 ( n17630 , n1852 , n17329 );
    or g10707 ( n19792 , n5277 , n2739 );
    not g10708 ( n26446 , n19979 );
    nor g10709 ( n15432 , n1802 , n18328 );
    not g10710 ( n12683 , n5038 );
    xnor g10711 ( n14054 , n3760 , n9860 );
    or g10712 ( n25055 , n2181 , n28866 );
    and g10713 ( n339 , n8429 , n11508 );
    or g10714 ( n16647 , n26388 , n22690 );
    or g10715 ( n2587 , n24066 , n23246 );
    or g10716 ( n31867 , n16839 , n8655 );
    xnor g10717 ( n14896 , n11413 , n4196 );
    or g10718 ( n7195 , n8998 , n9749 );
    xnor g10719 ( n19663 , n109 , n2001 );
    not g10720 ( n28222 , n17313 );
    xnor g10721 ( n15406 , n9580 , n9031 );
    or g10722 ( n20677 , n24709 , n18357 );
    nor g10723 ( n1011 , n23550 , n14463 );
    and g10724 ( n25638 , n22364 , n9936 );
    not g10725 ( n5045 , n3700 );
    not g10726 ( n25122 , n24198 );
    not g10727 ( n17854 , n4571 );
    and g10728 ( n25576 , n22198 , n12769 );
    buf g10729 ( n17917 , n29706 );
    and g10730 ( n29254 , n13409 , n26803 );
    xnor g10731 ( n17287 , n16410 , n1880 );
    xnor g10732 ( n2325 , n196 , n30930 );
    buf g10733 ( n4339 , n10019 );
    or g10734 ( n31399 , n26408 , n29282 );
    nor g10735 ( n16318 , n28036 , n27993 );
    and g10736 ( n20509 , n6706 , n16905 );
    or g10737 ( n17096 , n16109 , n31969 );
    xor g10738 ( n30453 , n27667 , n15929 );
    and g10739 ( n8000 , n4840 , n3266 );
    not g10740 ( n26507 , n21386 );
    xnor g10741 ( n23734 , n27804 , n945 );
    not g10742 ( n21879 , n28282 );
    or g10743 ( n27983 , n26009 , n15134 );
    not g10744 ( n3410 , n23750 );
    or g10745 ( n6567 , n3182 , n11906 );
    xnor g10746 ( n12435 , n20720 , n3510 );
    or g10747 ( n13557 , n1347 , n10504 );
    not g10748 ( n8334 , n2446 );
    or g10749 ( n38 , n3515 , n8300 );
    and g10750 ( n1814 , n7516 , n11275 );
    and g10751 ( n3539 , n13998 , n28397 );
    not g10752 ( n15401 , n5215 );
    xnor g10753 ( n2547 , n12836 , n2240 );
    or g10754 ( n27518 , n16495 , n15528 );
    nor g10755 ( n4104 , n13210 , n197 );
    xnor g10756 ( n19573 , n10850 , n16196 );
    nor g10757 ( n10918 , n29581 , n31323 );
    nor g10758 ( n9410 , n1997 , n12373 );
    not g10759 ( n14629 , n14361 );
    or g10760 ( n258 , n9582 , n17642 );
    not g10761 ( n30777 , n11781 );
    and g10762 ( n25565 , n21207 , n16743 );
    and g10763 ( n3136 , n9857 , n287 );
    or g10764 ( n21559 , n2470 , n24936 );
    or g10765 ( n10279 , n13367 , n21160 );
    or g10766 ( n18952 , n19140 , n18524 );
    nor g10767 ( n22165 , n19356 , n11423 );
    or g10768 ( n23808 , n24488 , n14829 );
    xnor g10769 ( n3270 , n20383 , n26381 );
    and g10770 ( n10999 , n27363 , n24952 );
    or g10771 ( n17323 , n19989 , n14650 );
    not g10772 ( n1040 , n7112 );
    or g10773 ( n26861 , n27746 , n18351 );
    xnor g10774 ( n324 , n16168 , n7775 );
    not g10775 ( n19982 , n23635 );
    not g10776 ( n29739 , n16468 );
    xor g10777 ( n20747 , n29225 , n24349 );
    not g10778 ( n30521 , n9070 );
    not g10779 ( n2613 , n19183 );
    nor g10780 ( n19210 , n26639 , n16942 );
    or g10781 ( n3041 , n20381 , n2708 );
    not g10782 ( n30380 , n6585 );
    xnor g10783 ( n7589 , n18042 , n5564 );
    or g10784 ( n27509 , n6196 , n5558 );
    not g10785 ( n5858 , n6692 );
    and g10786 ( n18358 , n5993 , n31282 );
    xnor g10787 ( n31206 , n25760 , n9239 );
    xnor g10788 ( n13400 , n28366 , n11039 );
    and g10789 ( n7348 , n26406 , n4994 );
    nor g10790 ( n11085 , n30486 , n27065 );
    not g10791 ( n15706 , n23252 );
    or g10792 ( n26282 , n428 , n26648 );
    xnor g10793 ( n15542 , n97 , n10451 );
    and g10794 ( n3205 , n5692 , n9534 );
    and g10795 ( n8534 , n10069 , n27243 );
    not g10796 ( n10707 , n2261 );
    or g10797 ( n4900 , n15793 , n25810 );
    and g10798 ( n23759 , n10318 , n4356 );
    not g10799 ( n15738 , n25774 );
    xnor g10800 ( n27433 , n24235 , n16441 );
    and g10801 ( n14192 , n1522 , n16744 );
    nor g10802 ( n8642 , n21597 , n19754 );
    or g10803 ( n27228 , n28824 , n23355 );
    xnor g10804 ( n11308 , n25863 , n1701 );
    or g10805 ( n9589 , n30297 , n1589 );
    or g10806 ( n24577 , n806 , n20479 );
    or g10807 ( n14809 , n23349 , n12451 );
    and g10808 ( n29979 , n12997 , n8674 );
    nor g10809 ( n24020 , n11792 , n27501 );
    and g10810 ( n19367 , n30452 , n20778 );
    not g10811 ( n5652 , n10165 );
    not g10812 ( n20657 , n16131 );
    and g10813 ( n6083 , n19214 , n30156 );
    xnor g10814 ( n16370 , n4231 , n6307 );
    or g10815 ( n13513 , n18891 , n17245 );
    not g10816 ( n30306 , n19951 );
    not g10817 ( n25843 , n14463 );
    not g10818 ( n25518 , n16254 );
    or g10819 ( n12408 , n12024 , n11671 );
    or g10820 ( n19461 , n7423 , n6560 );
    not g10821 ( n27916 , n23401 );
    and g10822 ( n24672 , n7439 , n23255 );
    not g10823 ( n2991 , n5250 );
    nor g10824 ( n28623 , n29659 , n21815 );
    and g10825 ( n912 , n11529 , n429 );
    not g10826 ( n8933 , n15531 );
    or g10827 ( n24623 , n25303 , n30077 );
    nor g10828 ( n24504 , n14230 , n23253 );
    or g10829 ( n28803 , n14133 , n20765 );
    and g10830 ( n16004 , n9252 , n22402 );
    not g10831 ( n27444 , n4836 );
    or g10832 ( n10470 , n4335 , n7559 );
    xnor g10833 ( n5732 , n1240 , n31999 );
    xnor g10834 ( n24531 , n15931 , n23382 );
    not g10835 ( n19368 , n27986 );
    not g10836 ( n5933 , n15125 );
    xnor g10837 ( n27272 , n25088 , n5475 );
    and g10838 ( n13589 , n27648 , n31713 );
    and g10839 ( n2298 , n19463 , n30252 );
    xnor g10840 ( n17333 , n935 , n21520 );
    or g10841 ( n1560 , n31562 , n1868 );
    or g10842 ( n31877 , n16603 , n5091 );
    or g10843 ( n7269 , n10427 , n2638 );
    not g10844 ( n14099 , n30808 );
    or g10845 ( n16377 , n28757 , n14637 );
    not g10846 ( n27484 , n5820 );
    or g10847 ( n16667 , n8753 , n18772 );
    nor g10848 ( n23755 , n16399 , n263 );
    not g10849 ( n27416 , n27925 );
    and g10850 ( n4613 , n1779 , n21045 );
    and g10851 ( n29971 , n2751 , n24741 );
    and g10852 ( n5899 , n19914 , n10940 );
    xnor g10853 ( n6217 , n16613 , n11430 );
    xnor g10854 ( n29285 , n18309 , n7683 );
    not g10855 ( n29100 , n8745 );
    and g10856 ( n18564 , n27421 , n5828 );
    nor g10857 ( n1564 , n5149 , n28297 );
    xnor g10858 ( n10929 , n30950 , n19738 );
    xnor g10859 ( n105 , n3714 , n9727 );
    xnor g10860 ( n8977 , n4268 , n11967 );
    or g10861 ( n8727 , n12663 , n14312 );
    xnor g10862 ( n20242 , n4007 , n29471 );
    not g10863 ( n30676 , n5646 );
    xnor g10864 ( n22037 , n12887 , n24525 );
    not g10865 ( n14128 , n26569 );
    or g10866 ( n30736 , n2898 , n12841 );
    xor g10867 ( n17835 , n30088 , n5402 );
    and g10868 ( n13195 , n1789 , n31167 );
    not g10869 ( n7194 , n12872 );
    xnor g10870 ( n8991 , n3499 , n9318 );
    or g10871 ( n28850 , n27590 , n1897 );
    xnor g10872 ( n14880 , n21991 , n6709 );
    or g10873 ( n11744 , n19429 , n26147 );
    nor g10874 ( n21288 , n21485 , n19373 );
    nor g10875 ( n3953 , n2135 , n18531 );
    or g10876 ( n14092 , n10984 , n21557 );
    xnor g10877 ( n28748 , n17777 , n25517 );
    not g10878 ( n5156 , n11393 );
    xnor g10879 ( n13488 , n5535 , n23578 );
    or g10880 ( n712 , n26548 , n28769 );
    xnor g10881 ( n1186 , n9638 , n13514 );
    buf g10882 ( n21272 , n12422 );
    not g10883 ( n15977 , n30381 );
    and g10884 ( n2479 , n29077 , n15123 );
    not g10885 ( n15311 , n4904 );
    xnor g10886 ( n30641 , n1267 , n29607 );
    not g10887 ( n8150 , n12075 );
    xnor g10888 ( n5166 , n27144 , n11658 );
    and g10889 ( n512 , n27561 , n16629 );
    xnor g10890 ( n17371 , n19513 , n24991 );
    or g10891 ( n23273 , n4275 , n362 );
    xnor g10892 ( n7600 , n7697 , n2347 );
    or g10893 ( n25951 , n5376 , n15969 );
    xnor g10894 ( n15763 , n26128 , n11735 );
    not g10895 ( n2315 , n4662 );
    and g10896 ( n29772 , n17725 , n12620 );
    or g10897 ( n28265 , n1370 , n20258 );
    nor g10898 ( n15129 , n27441 , n21902 );
    or g10899 ( n18680 , n25170 , n13565 );
    or g10900 ( n12599 , n10676 , n29745 );
    not g10901 ( n28867 , n29671 );
    xnor g10902 ( n28685 , n4287 , n2231 );
    not g10903 ( n22147 , n11543 );
    xnor g10904 ( n13276 , n13896 , n16403 );
    or g10905 ( n12539 , n19692 , n1418 );
    and g10906 ( n29213 , n14903 , n9227 );
    or g10907 ( n31161 , n12242 , n13999 );
    not g10908 ( n8491 , n3553 );
    not g10909 ( n22514 , n9485 );
    xnor g10910 ( n26292 , n11360 , n30067 );
    not g10911 ( n7677 , n19577 );
    and g10912 ( n3246 , n20571 , n21431 );
    or g10913 ( n16894 , n8987 , n5523 );
    xnor g10914 ( n1771 , n16132 , n891 );
    xnor g10915 ( n31672 , n13852 , n12946 );
    and g10916 ( n23593 , n18297 , n23656 );
    not g10917 ( n28297 , n16609 );
    xnor g10918 ( n10802 , n11184 , n26065 );
    not g10919 ( n3447 , n97 );
    or g10920 ( n14371 , n4946 , n20793 );
    xnor g10921 ( n27720 , n127 , n18007 );
    or g10922 ( n26042 , n28649 , n20915 );
    nor g10923 ( n10484 , n7525 , n21950 );
    and g10924 ( n24277 , n16243 , n6353 );
    xnor g10925 ( n26791 , n18645 , n18850 );
    not g10926 ( n19736 , n26173 );
    nor g10927 ( n14620 , n30684 , n612 );
    and g10928 ( n29055 , n13732 , n30519 );
    not g10929 ( n3597 , n22553 );
    or g10930 ( n186 , n5166 , n13503 );
    nor g10931 ( n12976 , n27432 , n26495 );
    and g10932 ( n13564 , n13605 , n18076 );
    or g10933 ( n27341 , n21824 , n6346 );
    xnor g10934 ( n13021 , n17282 , n28334 );
    or g10935 ( n9693 , n17481 , n28528 );
    xnor g10936 ( n9659 , n23735 , n13454 );
    and g10937 ( n13527 , n631 , n12539 );
    not g10938 ( n7360 , n7246 );
    not g10939 ( n13462 , n9040 );
    or g10940 ( n16680 , n6828 , n28396 );
    not g10941 ( n25319 , n1973 );
    xnor g10942 ( n25385 , n4616 , n24747 );
    or g10943 ( n889 , n8867 , n23777 );
    and g10944 ( n7665 , n331 , n29897 );
    or g10945 ( n361 , n28593 , n1410 );
    or g10946 ( n23038 , n3078 , n24966 );
    not g10947 ( n27084 , n3822 );
    and g10948 ( n20377 , n23501 , n16961 );
    or g10949 ( n8106 , n7241 , n29905 );
    and g10950 ( n24427 , n16691 , n26320 );
    not g10951 ( n20686 , n9642 );
    xnor g10952 ( n11845 , n30887 , n11771 );
    or g10953 ( n25663 , n26224 , n8516 );
    xnor g10954 ( n1170 , n22512 , n12668 );
    and g10955 ( n23923 , n15541 , n30834 );
    or g10956 ( n9252 , n24827 , n30701 );
    not g10957 ( n8613 , n5064 );
    or g10958 ( n16348 , n26966 , n19280 );
    not g10959 ( n25371 , n3169 );
    or g10960 ( n31314 , n7408 , n5847 );
    nor g10961 ( n9952 , n19006 , n28504 );
    not g10962 ( n15254 , n15854 );
    not g10963 ( n10716 , n27559 );
    and g10964 ( n16087 , n1684 , n14678 );
    and g10965 ( n21692 , n5462 , n23519 );
    and g10966 ( n16031 , n8583 , n24740 );
    and g10967 ( n5651 , n19528 , n19609 );
    xnor g10968 ( n3153 , n1050 , n10611 );
    nor g10969 ( n18802 , n11175 , n27831 );
    and g10970 ( n22468 , n6002 , n21384 );
    nor g10971 ( n8583 , n15823 , n17260 );
    xnor g10972 ( n21545 , n21797 , n15107 );
    not g10973 ( n29082 , n18538 );
    not g10974 ( n7672 , n20120 );
    not g10975 ( n15384 , n24583 );
    not g10976 ( n17475 , n25946 );
    and g10977 ( n26761 , n19650 , n29404 );
    and g10978 ( n2887 , n21211 , n12238 );
    not g10979 ( n3979 , n30340 );
    or g10980 ( n7975 , n18057 , n7487 );
    nor g10981 ( n20926 , n19405 , n16800 );
    and g10982 ( n30065 , n19049 , n11078 );
    nor g10983 ( n29889 , n14998 , n14787 );
    xnor g10984 ( n7771 , n28036 , n16843 );
    xnor g10985 ( n4117 , n3125 , n4471 );
    not g10986 ( n15755 , n11450 );
    and g10987 ( n32000 , n1820 , n27957 );
    not g10988 ( n28695 , n28923 );
    and g10989 ( n23632 , n28117 , n17142 );
    not g10990 ( n22157 , n31048 );
    and g10991 ( n6712 , n3037 , n30514 );
    or g10992 ( n14562 , n28094 , n9750 );
    or g10993 ( n20243 , n16815 , n27106 );
    not g10994 ( n2164 , n8017 );
    nor g10995 ( n19131 , n28012 , n13885 );
    not g10996 ( n17737 , n25007 );
    not g10997 ( n10538 , n4822 );
    xnor g10998 ( n5975 , n31358 , n17231 );
    xnor g10999 ( n4719 , n3398 , n5330 );
    xnor g11000 ( n3336 , n20379 , n27501 );
    xnor g11001 ( n17524 , n26045 , n4285 );
    or g11002 ( n29892 , n16408 , n23524 );
    xor g11003 ( n25235 , n10651 , n5227 );
    and g11004 ( n25368 , n5362 , n12797 );
    not g11005 ( n17095 , n18447 );
    or g11006 ( n18661 , n2183 , n6694 );
    xnor g11007 ( n20709 , n19641 , n25276 );
    not g11008 ( n28717 , n23614 );
    or g11009 ( n16159 , n1257 , n5253 );
    or g11010 ( n4078 , n29784 , n31159 );
    or g11011 ( n10940 , n18303 , n3429 );
    xnor g11012 ( n24829 , n1288 , n10934 );
    not g11013 ( n14892 , n14267 );
    or g11014 ( n21876 , n451 , n4571 );
    xnor g11015 ( n11284 , n25575 , n18515 );
    xnor g11016 ( n22564 , n16046 , n13958 );
    or g11017 ( n9316 , n14282 , n21164 );
    nor g11018 ( n29861 , n2453 , n7152 );
    and g11019 ( n3374 , n11678 , n17144 );
    not g11020 ( n19336 , n28512 );
    xnor g11021 ( n175 , n1285 , n30593 );
    xnor g11022 ( n26435 , n29197 , n21485 );
    xnor g11023 ( n19780 , n24552 , n22318 );
    not g11024 ( n1604 , n9424 );
    xnor g11025 ( n2846 , n14097 , n18624 );
    and g11026 ( n7244 , n17674 , n5979 );
    and g11027 ( n14706 , n7268 , n14878 );
    nor g11028 ( n10832 , n6315 , n17824 );
    or g11029 ( n20706 , n18388 , n17558 );
    xnor g11030 ( n17 , n8881 , n27514 );
    and g11031 ( n4105 , n7812 , n21087 );
    and g11032 ( n27878 , n22889 , n27280 );
    xnor g11033 ( n30544 , n14100 , n24132 );
    nor g11034 ( n31340 , n5578 , n22712 );
    not g11035 ( n3849 , n23699 );
    xnor g11036 ( n1246 , n22762 , n21950 );
    or g11037 ( n19781 , n9920 , n7282 );
    not g11038 ( n13493 , n5532 );
    and g11039 ( n411 , n22662 , n21361 );
    not g11040 ( n26592 , n22087 );
    or g11041 ( n4666 , n28991 , n3892 );
    xnor g11042 ( n30828 , n12579 , n367 );
    xnor g11043 ( n10370 , n24501 , n29445 );
    or g11044 ( n11827 , n7845 , n28761 );
    not g11045 ( n16397 , n17364 );
    not g11046 ( n11452 , n3934 );
    and g11047 ( n12358 , n16436 , n19238 );
    and g11048 ( n24027 , n28944 , n22880 );
    not g11049 ( n17661 , n26683 );
    not g11050 ( n31782 , n30664 );
    and g11051 ( n4884 , n12185 , n23298 );
    not g11052 ( n20190 , n16516 );
    xnor g11053 ( n22597 , n9396 , n17499 );
    or g11054 ( n15551 , n7434 , n14413 );
    or g11055 ( n29548 , n1923 , n30523 );
    not g11056 ( n7559 , n117 );
    or g11057 ( n6593 , n11386 , n4986 );
    not g11058 ( n24203 , n16848 );
    xnor g11059 ( n20715 , n3828 , n14504 );
    not g11060 ( n7427 , n24964 );
    or g11061 ( n24105 , n25082 , n14029 );
    and g11062 ( n18578 , n10346 , n12312 );
    not g11063 ( n15684 , n7655 );
    nor g11064 ( n8337 , n29175 , n6097 );
    xnor g11065 ( n11541 , n14328 , n9239 );
    nor g11066 ( n28645 , n7705 , n31111 );
    nor g11067 ( n19673 , n14124 , n2041 );
    xnor g11068 ( n14852 , n3515 , n16676 );
    and g11069 ( n24771 , n6272 , n25925 );
    not g11070 ( n10060 , n486 );
    xnor g11071 ( n8487 , n30139 , n25648 );
    xnor g11072 ( n16881 , n15455 , n24544 );
    and g11073 ( n12787 , n7268 , n16744 );
    or g11074 ( n10625 , n10270 , n6228 );
    not g11075 ( n3492 , n10466 );
    nor g11076 ( n7476 , n7651 , n11705 );
    nor g11077 ( n20993 , n11094 , n12898 );
    not g11078 ( n8802 , n20698 );
    and g11079 ( n18898 , n14215 , n5921 );
    and g11080 ( n17189 , n5804 , n3198 );
    not g11081 ( n27161 , n18893 );
    not g11082 ( n2216 , n2469 );
    not g11083 ( n6213 , n21875 );
    and g11084 ( n15227 , n19327 , n19578 );
    xnor g11085 ( n9484 , n17579 , n26002 );
    not g11086 ( n20472 , n26271 );
    not g11087 ( n6061 , n15526 );
    or g11088 ( n22670 , n21935 , n6982 );
    nor g11089 ( n10526 , n31972 , n16930 );
    and g11090 ( n4420 , n27007 , n28316 );
    and g11091 ( n5841 , n12939 , n9900 );
    not g11092 ( n3920 , n26690 );
    and g11093 ( n77 , n6846 , n6693 );
    not g11094 ( n21172 , n25278 );
    nor g11095 ( n11989 , n19516 , n3299 );
    or g11096 ( n24310 , n8965 , n28478 );
    xnor g11097 ( n31450 , n15861 , n17910 );
    not g11098 ( n10776 , n23058 );
    nor g11099 ( n30456 , n21025 , n21723 );
    or g11100 ( n22783 , n1428 , n15243 );
    not g11101 ( n31085 , n23757 );
    not g11102 ( n21085 , n24750 );
    and g11103 ( n22463 , n8366 , n21766 );
    or g11104 ( n30708 , n12813 , n23584 );
    or g11105 ( n22038 , n21458 , n3926 );
    and g11106 ( n557 , n9420 , n18223 );
    xnor g11107 ( n30742 , n20574 , n1146 );
    or g11108 ( n28452 , n143 , n16628 );
    xnor g11109 ( n18589 , n27434 , n4844 );
    not g11110 ( n18548 , n26306 );
    nor g11111 ( n13304 , n7006 , n22046 );
    or g11112 ( n20533 , n13635 , n3929 );
    or g11113 ( n8674 , n16625 , n3171 );
    nor g11114 ( n18024 , n21523 , n6483 );
    or g11115 ( n0 , n26028 , n21238 );
    buf g11116 ( n5715 , n5125 );
    not g11117 ( n12016 , n7709 );
    xnor g11118 ( n26068 , n28566 , n9340 );
    not g11119 ( n27037 , n11692 );
    and g11120 ( n6055 , n10608 , n24437 );
    not g11121 ( n13429 , n27979 );
    nor g11122 ( n13401 , n22917 , n3345 );
    xnor g11123 ( n23353 , n5477 , n4665 );
    xnor g11124 ( n30113 , n17008 , n24063 );
    and g11125 ( n2768 , n3520 , n9570 );
    and g11126 ( n9330 , n30194 , n7318 );
    not g11127 ( n27821 , n1031 );
    not g11128 ( n15563 , n23561 );
    xnor g11129 ( n23941 , n30864 , n11527 );
    or g11130 ( n15600 , n21485 , n6488 );
    not g11131 ( n25481 , n30911 );
    nor g11132 ( n29177 , n6121 , n7248 );
    and g11133 ( n18664 , n15462 , n13413 );
    or g11134 ( n30140 , n16183 , n15679 );
    xnor g11135 ( n23323 , n933 , n20667 );
    xnor g11136 ( n19149 , n12606 , n14163 );
    and g11137 ( n3237 , n28876 , n4293 );
    xnor g11138 ( n29458 , n9744 , n15382 );
    xnor g11139 ( n4708 , n19760 , n30181 );
    not g11140 ( n28050 , n12941 );
    and g11141 ( n3477 , n8650 , n1556 );
    not g11142 ( n9912 , n9071 );
    not g11143 ( n7022 , n3613 );
    xnor g11144 ( n28943 , n21811 , n31173 );
    or g11145 ( n1189 , n30117 , n23951 );
    xor g11146 ( n9472 , n17121 , n8093 );
    not g11147 ( n10747 , n25444 );
    and g11148 ( n14125 , n11589 , n21894 );
    nor g11149 ( n3271 , n13318 , n28159 );
    and g11150 ( n13189 , n12890 , n15147 );
    and g11151 ( n25655 , n31706 , n8859 );
    nor g11152 ( n465 , n8234 , n16541 );
    not g11153 ( n1698 , n9660 );
    xnor g11154 ( n4630 , n27693 , n27077 );
    xnor g11155 ( n28953 , n30244 , n19007 );
    not g11156 ( n26762 , n14269 );
    not g11157 ( n15514 , n17966 );
    xnor g11158 ( n10690 , n12228 , n19676 );
    xnor g11159 ( n182 , n16486 , n17726 );
    and g11160 ( n11501 , n18205 , n16611 );
    or g11161 ( n6299 , n6989 , n7273 );
    and g11162 ( n3055 , n29613 , n23000 );
    nor g11163 ( n13853 , n28081 , n785 );
    not g11164 ( n11709 , n15797 );
    not g11165 ( n6695 , n30071 );
    not g11166 ( n2180 , n9612 );
    or g11167 ( n16130 , n1970 , n28304 );
    and g11168 ( n3972 , n5829 , n12748 );
    not g11169 ( n23129 , n4458 );
    or g11170 ( n13033 , n13860 , n30403 );
    not g11171 ( n12053 , n5684 );
    or g11172 ( n4234 , n13979 , n23805 );
    and g11173 ( n20794 , n24945 , n22334 );
    or g11174 ( n10231 , n3065 , n19743 );
    or g11175 ( n18386 , n3676 , n9351 );
    or g11176 ( n7106 , n30165 , n8434 );
    or g11177 ( n17011 , n11436 , n21328 );
    or g11178 ( n16502 , n5685 , n6968 );
    not g11179 ( n2998 , n30695 );
    xnor g11180 ( n27015 , n18327 , n2883 );
    xnor g11181 ( n26123 , n30067 , n9338 );
    and g11182 ( n26140 , n15268 , n28411 );
    and g11183 ( n12904 , n14022 , n27158 );
    or g11184 ( n3026 , n26536 , n10187 );
    xnor g11185 ( n20296 , n21136 , n31366 );
    not g11186 ( n9586 , n30775 );
    xnor g11187 ( n851 , n4456 , n25291 );
    or g11188 ( n30844 , n25425 , n10982 );
    and g11189 ( n28701 , n20935 , n27488 );
    and g11190 ( n8661 , n839 , n13143 );
    xnor g11191 ( n2262 , n16862 , n13975 );
    not g11192 ( n11280 , n22817 );
    xnor g11193 ( n23281 , n24132 , n29897 );
    and g11194 ( n15633 , n21769 , n28075 );
    not g11195 ( n4246 , n24118 );
    not g11196 ( n13930 , n3991 );
    nor g11197 ( n23911 , n30048 , n4650 );
    or g11198 ( n15656 , n27018 , n29856 );
    xnor g11199 ( n1987 , n11500 , n2126 );
    or g11200 ( n23105 , n20267 , n13354 );
    not g11201 ( n21463 , n15091 );
    or g11202 ( n28074 , n15187 , n1824 );
    not g11203 ( n12052 , n13877 );
    nor g11204 ( n1991 , n10269 , n17248 );
    nor g11205 ( n31850 , n30313 , n30578 );
    xnor g11206 ( n23936 , n3080 , n2934 );
    nor g11207 ( n13941 , n29759 , n18688 );
    or g11208 ( n31356 , n19130 , n8209 );
    nor g11209 ( n30700 , n30014 , n15334 );
    or g11210 ( n15005 , n15172 , n12367 );
    or g11211 ( n16018 , n864 , n10828 );
    not g11212 ( n26491 , n31707 );
    xnor g11213 ( n9535 , n7416 , n30502 );
    not g11214 ( n9047 , n29854 );
    or g11215 ( n17120 , n8826 , n7497 );
    and g11216 ( n27969 , n11053 , n24424 );
    not g11217 ( n2727 , n13003 );
    xnor g11218 ( n31267 , n316 , n8987 );
    not g11219 ( n7621 , n26481 );
    and g11220 ( n10572 , n3918 , n30539 );
    not g11221 ( n6965 , n7208 );
    and g11222 ( n22158 , n5091 , n16603 );
    or g11223 ( n24270 , n23160 , n23483 );
    not g11224 ( n4684 , n12412 );
    not g11225 ( n22245 , n14015 );
    not g11226 ( n21678 , n8872 );
    and g11227 ( n30422 , n20883 , n8901 );
    or g11228 ( n5224 , n31318 , n14743 );
    nor g11229 ( n28656 , n14026 , n17131 );
    xnor g11230 ( n28374 , n21900 , n23538 );
    xnor g11231 ( n5297 , n3131 , n20881 );
    not g11232 ( n5747 , n26592 );
    or g11233 ( n464 , n31111 , n27067 );
    xnor g11234 ( n11230 , n10573 , n9634 );
    xnor g11235 ( n14380 , n13198 , n19746 );
    nor g11236 ( n19628 , n27077 , n12207 );
    xnor g11237 ( n19354 , n8767 , n4710 );
    or g11238 ( n26372 , n9623 , n29240 );
    xnor g11239 ( n5560 , n13482 , n9975 );
    not g11240 ( n12183 , n28579 );
    and g11241 ( n5626 , n10328 , n23136 );
    not g11242 ( n8098 , n8338 );
    xnor g11243 ( n17342 , n26116 , n19788 );
    not g11244 ( n17842 , n3943 );
    not g11245 ( n31128 , n27529 );
    buf g11246 ( n209 , n12199 );
    nor g11247 ( n21060 , n3752 , n12866 );
    xnor g11248 ( n19852 , n22068 , n14277 );
    not g11249 ( n21841 , n2339 );
    not g11250 ( n17253 , n5092 );
    xnor g11251 ( n14208 , n26683 , n5974 );
    or g11252 ( n4880 , n17703 , n30527 );
    and g11253 ( n9117 , n31530 , n8448 );
    and g11254 ( n19304 , n13600 , n30356 );
    and g11255 ( n30170 , n8182 , n5291 );
    nor g11256 ( n9072 , n14925 , n25393 );
    not g11257 ( n18210 , n5831 );
    xnor g11258 ( n21391 , n22233 , n25760 );
    not g11259 ( n23182 , n25660 );
    or g11260 ( n28893 , n19079 , n16188 );
    buf g11261 ( n24225 , n19094 );
    and g11262 ( n22578 , n669 , n10334 );
    xnor g11263 ( n2804 , n15199 , n26807 );
    xnor g11264 ( n16192 , n3543 , n1458 );
    or g11265 ( n2497 , n3840 , n29204 );
    not g11266 ( n18017 , n85 );
    or g11267 ( n30100 , n1412 , n22728 );
    not g11268 ( n30029 , n13560 );
    and g11269 ( n9250 , n15094 , n3022 );
    nor g11270 ( n11881 , n25454 , n4074 );
    not g11271 ( n13326 , n876 );
    not g11272 ( n6998 , n9310 );
    nor g11273 ( n28780 , n18778 , n30917 );
    nor g11274 ( n4141 , n5387 , n6295 );
    and g11275 ( n5796 , n31664 , n21603 );
    not g11276 ( n21638 , n11721 );
    not g11277 ( n8388 , n12346 );
    xnor g11278 ( n17715 , n24396 , n21023 );
    buf g11279 ( n674 , n14610 );
    not g11280 ( n11057 , n8672 );
    or g11281 ( n8788 , n11314 , n30400 );
    xnor g11282 ( n739 , n25885 , n14929 );
    and g11283 ( n3855 , n9020 , n1200 );
    xnor g11284 ( n15802 , n30961 , n8934 );
    nor g11285 ( n18145 , n2753 , n8311 );
    or g11286 ( n191 , n30386 , n20294 );
    xor g11287 ( n2588 , n1929 , n19548 );
    xnor g11288 ( n27129 , n31786 , n8901 );
    xnor g11289 ( n7749 , n2910 , n16406 );
    xnor g11290 ( n1272 , n3036 , n26004 );
    or g11291 ( n2133 , n14076 , n13706 );
    or g11292 ( n19473 , n30601 , n8562 );
    or g11293 ( n17583 , n8331 , n19876 );
    or g11294 ( n20585 , n13494 , n30519 );
    nor g11295 ( n17240 , n27152 , n26343 );
    not g11296 ( n9383 , n8346 );
    xnor g11297 ( n14591 , n10123 , n807 );
    not g11298 ( n4128 , n9572 );
    xnor g11299 ( n6427 , n22404 , n10190 );
    and g11300 ( n17494 , n14855 , n5537 );
    and g11301 ( n8212 , n22353 , n17258 );
    or g11302 ( n3104 , n27534 , n10981 );
    xnor g11303 ( n29986 , n22870 , n2444 );
    not g11304 ( n700 , n26495 );
    not g11305 ( n6361 , n5608 );
    and g11306 ( n29957 , n25787 , n4063 );
    and g11307 ( n2203 , n11922 , n8192 );
    and g11308 ( n29625 , n22638 , n25956 );
    and g11309 ( n14261 , n22026 , n27297 );
    or g11310 ( n18277 , n8260 , n31905 );
    not g11311 ( n15321 , n20982 );
    or g11312 ( n1553 , n24687 , n4134 );
    nor g11313 ( n10313 , n19500 , n28665 );
    not g11314 ( n3195 , n515 );
    and g11315 ( n23352 , n16035 , n12517 );
    and g11316 ( n3667 , n25118 , n7786 );
    and g11317 ( n7186 , n14909 , n4391 );
    not g11318 ( n30270 , n17981 );
    and g11319 ( n376 , n10811 , n24434 );
    or g11320 ( n6281 , n10283 , n10675 );
    not g11321 ( n9177 , n31353 );
    or g11322 ( n10784 , n23070 , n17752 );
    xnor g11323 ( n21787 , n7462 , n30735 );
    xor g11324 ( n13235 , n10234 , n7743 );
    nor g11325 ( n1511 , n30769 , n9312 );
    xnor g11326 ( n3096 , n12096 , n16193 );
    or g11327 ( n11556 , n26419 , n3866 );
    or g11328 ( n10349 , n7861 , n11700 );
    and g11329 ( n16613 , n10968 , n1735 );
    xnor g11330 ( n2300 , n10071 , n9835 );
    xor g11331 ( n17150 , n16746 , n28758 );
    not g11332 ( n8071 , n8413 );
    nor g11333 ( n17208 , n28828 , n6196 );
    or g11334 ( n25830 , n26867 , n16958 );
    and g11335 ( n26340 , n18607 , n8262 );
    xnor g11336 ( n1062 , n11030 , n12601 );
    xnor g11337 ( n14421 , n18154 , n22863 );
    or g11338 ( n17967 , n19247 , n4731 );
    or g11339 ( n21236 , n7356 , n28099 );
    not g11340 ( n2143 , n2105 );
    or g11341 ( n15537 , n1770 , n2291 );
    and g11342 ( n10065 , n5667 , n11249 );
    not g11343 ( n8357 , n2291 );
    or g11344 ( n9511 , n12624 , n9333 );
    or g11345 ( n6847 , n23116 , n21112 );
    or g11346 ( n7296 , n14927 , n3874 );
    not g11347 ( n16747 , n12340 );
    xnor g11348 ( n1146 , n11842 , n14141 );
    nor g11349 ( n20413 , n2855 , n12147 );
    or g11350 ( n30559 , n15399 , n28563 );
    or g11351 ( n5021 , n15624 , n22522 );
    nor g11352 ( n22825 , n13454 , n13724 );
    not g11353 ( n2990 , n2461 );
    not g11354 ( n29483 , n9031 );
    xnor g11355 ( n24114 , n1469 , n29037 );
    not g11356 ( n29527 , n28531 );
    not g11357 ( n23889 , n15439 );
    and g11358 ( n637 , n3677 , n24481 );
    and g11359 ( n28097 , n7441 , n25411 );
    and g11360 ( n17861 , n26345 , n24615 );
    not g11361 ( n2188 , n17772 );
    nor g11362 ( n16082 , n26409 , n23608 );
    not g11363 ( n10208 , n3160 );
    or g11364 ( n20681 , n1366 , n4439 );
    not g11365 ( n16360 , n27632 );
    and g11366 ( n20991 , n2927 , n1362 );
    xnor g11367 ( n15152 , n21559 , n3781 );
    xnor g11368 ( n6628 , n11220 , n32024 );
    nor g11369 ( n11787 , n26313 , n1173 );
    not g11370 ( n25677 , n26052 );
    nor g11371 ( n27229 , n11026 , n15113 );
    or g11372 ( n24281 , n25298 , n28721 );
    xnor g11373 ( n2336 , n30777 , n25334 );
    not g11374 ( n6599 , n6489 );
    or g11375 ( n28650 , n19122 , n1627 );
    nor g11376 ( n30118 , n30535 , n26620 );
    nor g11377 ( n2554 , n5779 , n13666 );
    and g11378 ( n2607 , n9523 , n14757 );
    not g11379 ( n2169 , n14387 );
    not g11380 ( n792 , n8778 );
    or g11381 ( n8621 , n29786 , n25071 );
    xnor g11382 ( n24892 , n5507 , n13355 );
    xnor g11383 ( n9202 , n216 , n18727 );
    or g11384 ( n27212 , n13226 , n23993 );
    xnor g11385 ( n28681 , n8184 , n2398 );
    not g11386 ( n29845 , n7240 );
    not g11387 ( n3914 , n9832 );
    and g11388 ( n28933 , n13253 , n17660 );
    or g11389 ( n25068 , n15673 , n27290 );
    xnor g11390 ( n16471 , n20826 , n2799 );
    buf g11391 ( n30045 , n30186 );
    or g11392 ( n24763 , n14199 , n29383 );
    or g11393 ( n7556 , n11420 , n5106 );
    or g11394 ( n17400 , n15700 , n8065 );
    xnor g11395 ( n1251 , n23071 , n18516 );
    or g11396 ( n7364 , n27779 , n5891 );
    xnor g11397 ( n5884 , n17478 , n3584 );
    not g11398 ( n9401 , n7351 );
    not g11399 ( n16934 , n6610 );
    xnor g11400 ( n20144 , n15716 , n23256 );
    or g11401 ( n24677 , n22571 , n14516 );
    or g11402 ( n17273 , n24498 , n7312 );
    xnor g11403 ( n28604 , n16606 , n15274 );
    xnor g11404 ( n27970 , n22867 , n12030 );
    not g11405 ( n9219 , n8991 );
    and g11406 ( n17256 , n18306 , n5623 );
    or g11407 ( n22797 , n22161 , n27209 );
    xnor g11408 ( n29671 , n2733 , n3331 );
    not g11409 ( n25425 , n24687 );
    not g11410 ( n27796 , n11826 );
    xnor g11411 ( n27206 , n1616 , n21597 );
    xor g11412 ( n20480 , n639 , n20446 );
    xor g11413 ( n3624 , n14321 , n15998 );
    nor g11414 ( n19809 , n25832 , n19067 );
    xnor g11415 ( n6707 , n14833 , n14609 );
    not g11416 ( n19033 , n1977 );
    not g11417 ( n28492 , n14441 );
    or g11418 ( n10459 , n5471 , n4339 );
    not g11419 ( n2856 , n15111 );
    not g11420 ( n27574 , n1012 );
    not g11421 ( n28010 , n28437 );
    not g11422 ( n13296 , n13147 );
    not g11423 ( n28440 , n29249 );
    nor g11424 ( n27645 , n22512 , n16956 );
    xnor g11425 ( n7766 , n3782 , n27354 );
    not g11426 ( n25581 , n1430 );
    and g11427 ( n7887 , n6461 , n22038 );
    not g11428 ( n13897 , n14999 );
    nor g11429 ( n21761 , n20438 , n203 );
    or g11430 ( n14478 , n31169 , n30928 );
    not g11431 ( n28302 , n4854 );
    xnor g11432 ( n4703 , n15778 , n1635 );
    xnor g11433 ( n348 , n1657 , n31765 );
    or g11434 ( n26753 , n14577 , n8290 );
    xnor g11435 ( n9880 , n25876 , n2325 );
    not g11436 ( n10483 , n10638 );
    not g11437 ( n25648 , n12407 );
    or g11438 ( n8652 , n15993 , n20113 );
    and g11439 ( n26776 , n15319 , n19064 );
    nor g11440 ( n4492 , n28417 , n15252 );
    not g11441 ( n6923 , n7637 );
    xnor g11442 ( n16124 , n19583 , n27951 );
    not g11443 ( n21099 , n30856 );
    nor g11444 ( n17602 , n10982 , n31303 );
    or g11445 ( n22327 , n17886 , n22832 );
    xnor g11446 ( n27455 , n2897 , n30448 );
    xor g11447 ( n2370 , n19009 , n3252 );
    or g11448 ( n14486 , n21869 , n14558 );
    not g11449 ( n19434 , n461 );
    xnor g11450 ( n25199 , n10291 , n20240 );
    xnor g11451 ( n683 , n3226 , n27806 );
    and g11452 ( n7696 , n2668 , n7552 );
    and g11453 ( n10009 , n25022 , n4797 );
    not g11454 ( n17654 , n2751 );
    not g11455 ( n11246 , n22857 );
    or g11456 ( n12996 , n14720 , n2388 );
    nor g11457 ( n15935 , n238 , n28413 );
    and g11458 ( n24483 , n24454 , n2096 );
    or g11459 ( n14730 , n6556 , n1303 );
    not g11460 ( n24776 , n22496 );
    not g11461 ( n23520 , n18211 );
    xnor g11462 ( n19099 , n24487 , n7692 );
    xor g11463 ( n24827 , n4535 , n25234 );
    nor g11464 ( n3977 , n29426 , n2682 );
    or g11465 ( n26838 , n24400 , n4814 );
    nor g11466 ( n22133 , n31448 , n11984 );
    not g11467 ( n16810 , n19311 );
    and g11468 ( n18868 , n31089 , n20928 );
    not g11469 ( n5386 , n10933 );
    or g11470 ( n2500 , n28134 , n21781 );
    not g11471 ( n12151 , n19014 );
    xnor g11472 ( n19591 , n7402 , n29901 );
    xnor g11473 ( n927 , n20081 , n19610 );
    or g11474 ( n31547 , n7256 , n14978 );
    not g11475 ( n13659 , n24675 );
    xnor g11476 ( n12073 , n6724 , n232 );
    xnor g11477 ( n16090 , n15987 , n30514 );
    not g11478 ( n15073 , n20804 );
    not g11479 ( n22339 , n28611 );
    not g11480 ( n1994 , n13083 );
    nor g11481 ( n14890 , n22746 , n31489 );
    not g11482 ( n24057 , n11966 );
    nor g11483 ( n3444 , n26006 , n7017 );
    or g11484 ( n18844 , n4129 , n17680 );
    not g11485 ( n8512 , n29966 );
    not g11486 ( n31188 , n28896 );
    or g11487 ( n7936 , n6266 , n5818 );
    and g11488 ( n6186 , n12164 , n26685 );
    and g11489 ( n8040 , n20087 , n12309 );
    not g11490 ( n15159 , n30568 );
    nor g11491 ( n22724 , n1039 , n23024 );
    not g11492 ( n22103 , n23381 );
    and g11493 ( n29856 , n2619 , n17204 );
    xnor g11494 ( n26595 , n10818 , n7219 );
    and g11495 ( n11872 , n21118 , n47 );
    xnor g11496 ( n9058 , n18724 , n11701 );
    or g11497 ( n25302 , n5618 , n22272 );
    or g11498 ( n7853 , n31620 , n9048 );
    or g11499 ( n5832 , n17289 , n8359 );
    xnor g11500 ( n16454 , n14513 , n181 );
    not g11501 ( n20108 , n23019 );
    xnor g11502 ( n12601 , n14986 , n15760 );
    xnor g11503 ( n2655 , n5391 , n13332 );
    and g11504 ( n30316 , n16297 , n2504 );
    not g11505 ( n25547 , n1040 );
    xnor g11506 ( n26987 , n9763 , n20905 );
    nor g11507 ( n13047 , n26191 , n17910 );
    xnor g11508 ( n15578 , n16867 , n1856 );
    not g11509 ( n19160 , n21253 );
    and g11510 ( n2850 , n14893 , n9403 );
    nor g11511 ( n11404 , n28194 , n10944 );
    xnor g11512 ( n28451 , n13609 , n31372 );
    not g11513 ( n27326 , n11494 );
    not g11514 ( n19078 , n18452 );
    not g11515 ( n23368 , n23218 );
    nor g11516 ( n7713 , n11551 , n28162 );
    nor g11517 ( n6048 , n3858 , n20116 );
    or g11518 ( n4162 , n8342 , n6622 );
    xnor g11519 ( n23389 , n28359 , n11970 );
    xnor g11520 ( n31000 , n136 , n22471 );
    nor g11521 ( n12113 , n9948 , n9396 );
    or g11522 ( n15994 , n23306 , n9935 );
    not g11523 ( n21210 , n4847 );
    not g11524 ( n1296 , n28816 );
    not g11525 ( n15332 , n7778 );
    or g11526 ( n21978 , n15706 , n23931 );
    xnor g11527 ( n6133 , n28941 , n21234 );
    and g11528 ( n7060 , n26816 , n27465 );
    xnor g11529 ( n10610 , n4623 , n20453 );
    and g11530 ( n12415 , n17129 , n8643 );
    buf g11531 ( n11305 , n6610 );
    or g11532 ( n7305 , n19176 , n13792 );
    xnor g11533 ( n25150 , n335 , n9146 );
    and g11534 ( n1419 , n6674 , n350 );
    xnor g11535 ( n20295 , n23247 , n1683 );
    nor g11536 ( n31342 , n30287 , n9336 );
    nor g11537 ( n4609 , n19255 , n27444 );
    not g11538 ( n21259 , n25333 );
    or g11539 ( n11955 , n10421 , n6457 );
    nor g11540 ( n25841 , n23921 , n27481 );
    nor g11541 ( n30584 , n21743 , n18681 );
    and g11542 ( n12114 , n23168 , n4806 );
    xnor g11543 ( n8208 , n3297 , n9619 );
    or g11544 ( n17838 , n18409 , n15019 );
    and g11545 ( n11397 , n11190 , n31531 );
    not g11546 ( n21925 , n300 );
    xor g11547 ( n17441 , n2622 , n8559 );
    xnor g11548 ( n24593 , n22738 , n8713 );
    not g11549 ( n2241 , n25064 );
    xnor g11550 ( n28552 , n9761 , n17780 );
    or g11551 ( n22337 , n29085 , n26340 );
    nor g11552 ( n19931 , n3810 , n1479 );
    or g11553 ( n7490 , n27303 , n8050 );
    or g11554 ( n23930 , n30924 , n17681 );
    not g11555 ( n28914 , n9938 );
    xnor g11556 ( n11402 , n11125 , n19233 );
    not g11557 ( n23249 , n17306 );
    or g11558 ( n8174 , n11414 , n3939 );
    not g11559 ( n18886 , n20916 );
    xnor g11560 ( n12231 , n8717 , n23885 );
    or g11561 ( n24233 , n14475 , n30045 );
    not g11562 ( n312 , n10497 );
    not g11563 ( n27043 , n17969 );
    xnor g11564 ( n27010 , n27929 , n31076 );
    and g11565 ( n8805 , n9004 , n20851 );
    and g11566 ( n12173 , n16029 , n2555 );
    xnor g11567 ( n21358 , n10666 , n10529 );
    xnor g11568 ( n2964 , n22512 , n6874 );
    nor g11569 ( n15883 , n26961 , n2026 );
    xnor g11570 ( n16431 , n31112 , n20160 );
    xnor g11571 ( n8296 , n8044 , n30169 );
    xnor g11572 ( n4728 , n29892 , n19170 );
    and g11573 ( n30765 , n10533 , n7110 );
    or g11574 ( n9957 , n21078 , n31245 );
    not g11575 ( n1414 , n14385 );
    xor g11576 ( n13568 , n16842 , n29087 );
    and g11577 ( n20802 , n30926 , n15590 );
    not g11578 ( n31651 , n30273 );
    nor g11579 ( n5621 , n18972 , n23626 );
    or g11580 ( n9869 , n27980 , n13630 );
    xnor g11581 ( n18623 , n30966 , n9944 );
    or g11582 ( n7443 , n14377 , n29237 );
    xnor g11583 ( n8791 , n28690 , n21223 );
    or g11584 ( n25751 , n27610 , n20868 );
    not g11585 ( n29678 , n21525 );
    not g11586 ( n4897 , n20176 );
    not g11587 ( n11421 , n6704 );
    xnor g11588 ( n4026 , n28217 , n31156 );
    and g11589 ( n27099 , n25640 , n2561 );
    xnor g11590 ( n2652 , n14278 , n15501 );
    nor g11591 ( n25482 , n7855 , n4739 );
    or g11592 ( n19894 , n25589 , n1207 );
    xnor g11593 ( n12092 , n27355 , n24525 );
    nor g11594 ( n93 , n1433 , n29116 );
    not g11595 ( n9739 , n20031 );
    or g11596 ( n25822 , n20059 , n16097 );
    not g11597 ( n19536 , n4248 );
    xnor g11598 ( n13278 , n11736 , n5873 );
    and g11599 ( n6122 , n2241 , n1093 );
    or g11600 ( n12923 , n13407 , n29213 );
    xnor g11601 ( n30028 , n30906 , n4213 );
    xnor g11602 ( n29194 , n7452 , n11047 );
    not g11603 ( n20460 , n22065 );
    xnor g11604 ( n27928 , n19956 , n9831 );
    or g11605 ( n12295 , n25758 , n30292 );
    xnor g11606 ( n13887 , n3012 , n17992 );
    and g11607 ( n5966 , n27784 , n17981 );
    nor g11608 ( n18295 , n29834 , n3626 );
    nor g11609 ( n11142 , n30425 , n6243 );
    or g11610 ( n8304 , n11125 , n4637 );
    not g11611 ( n2634 , n4734 );
    nor g11612 ( n22749 , n4957 , n31363 );
    xnor g11613 ( n21870 , n28698 , n4863 );
    or g11614 ( n20419 , n17888 , n10561 );
    not g11615 ( n13857 , n29083 );
    xnor g11616 ( n9370 , n15393 , n29718 );
    not g11617 ( n2681 , n5288 );
    not g11618 ( n16689 , n3822 );
    or g11619 ( n29698 , n932 , n28192 );
    nor g11620 ( n10198 , n20538 , n274 );
    and g11621 ( n5121 , n14660 , n3521 );
    not g11622 ( n13171 , n30037 );
    xnor g11623 ( n3228 , n13532 , n23353 );
    not g11624 ( n5339 , n25699 );
    or g11625 ( n3891 , n6832 , n9644 );
    not g11626 ( n14923 , n12169 );
    or g11627 ( n31774 , n4391 , n21379 );
    nor g11628 ( n8291 , n25262 , n24993 );
    not g11629 ( n22156 , n11610 );
    xnor g11630 ( n16101 , n22997 , n14025 );
    not g11631 ( n2021 , n9141 );
    and g11632 ( n13909 , n30598 , n7678 );
    or g11633 ( n26847 , n25218 , n11965 );
    not g11634 ( n12169 , n4968 );
    not g11635 ( n3861 , n27176 );
    and g11636 ( n16263 , n21069 , n12735 );
    xnor g11637 ( n677 , n30638 , n20844 );
    and g11638 ( n24919 , n30372 , n7609 );
    or g11639 ( n24252 , n10373 , n28143 );
    nor g11640 ( n16439 , n12929 , n31216 );
    xnor g11641 ( n15976 , n30412 , n11197 );
    buf g11642 ( n17166 , n20980 );
    or g11643 ( n19163 , n17467 , n2735 );
    xnor g11644 ( n4254 , n18004 , n19182 );
    not g11645 ( n28036 , n13260 );
    not g11646 ( n2625 , n16406 );
    and g11647 ( n29149 , n21052 , n2892 );
    and g11648 ( n5408 , n26397 , n27900 );
    not g11649 ( n28715 , n17115 );
    and g11650 ( n14006 , n7615 , n21451 );
    not g11651 ( n26100 , n3832 );
    xnor g11652 ( n29001 , n18310 , n5884 );
    nor g11653 ( n16880 , n17158 , n26688 );
    or g11654 ( n3732 , n22538 , n3260 );
    or g11655 ( n16976 , n12013 , n2131 );
    not g11656 ( n101 , n23974 );
    or g11657 ( n10265 , n3603 , n22103 );
    not g11658 ( n6115 , n6199 );
    or g11659 ( n1655 , n10822 , n2436 );
    not g11660 ( n1956 , n2236 );
    xnor g11661 ( n18657 , n13063 , n18394 );
    and g11662 ( n31859 , n18222 , n24073 );
    or g11663 ( n5645 , n21579 , n4445 );
    not g11664 ( n20218 , n27062 );
    nor g11665 ( n26677 , n26786 , n11799 );
    not g11666 ( n16581 , n22549 );
    not g11667 ( n2844 , n3854 );
    xnor g11668 ( n26579 , n9407 , n7825 );
    and g11669 ( n22507 , n24293 , n6625 );
    xor g11670 ( n19177 , n11959 , n26289 );
    and g11671 ( n2048 , n9321 , n26863 );
    xnor g11672 ( n18003 , n13503 , n6327 );
    xnor g11673 ( n24999 , n3107 , n18140 );
    not g11674 ( n26901 , n26162 );
    not g11675 ( n5826 , n607 );
    or g11676 ( n25916 , n14416 , n4181 );
    buf g11677 ( n5924 , n6082 );
    not g11678 ( n3154 , n6554 );
    not g11679 ( n7127 , n26082 );
    not g11680 ( n14942 , n16288 );
    xnor g11681 ( n29967 , n13202 , n5766 );
    not g11682 ( n28851 , n22434 );
    or g11683 ( n13637 , n16861 , n28532 );
    or g11684 ( n30531 , n24464 , n2410 );
    or g11685 ( n18212 , n28983 , n30014 );
    and g11686 ( n12536 , n9884 , n9934 );
    or g11687 ( n27082 , n3975 , n22087 );
    xor g11688 ( n31386 , n29246 , n30296 );
    or g11689 ( n9161 , n28441 , n21621 );
    xnor g11690 ( n11634 , n2479 , n22871 );
    xnor g11691 ( n27056 , n3603 , n27088 );
    xnor g11692 ( n6505 , n15343 , n23979 );
    xnor g11693 ( n23997 , n18906 , n29072 );
    xnor g11694 ( n2726 , n25558 , n16998 );
    and g11695 ( n31035 , n6917 , n28238 );
    not g11696 ( n30184 , n25562 );
    not g11697 ( n7124 , n1388 );
    and g11698 ( n17549 , n8375 , n26701 );
    and g11699 ( n14031 , n22050 , n14746 );
    not g11700 ( n27221 , n22434 );
    or g11701 ( n7811 , n12439 , n30958 );
    xnor g11702 ( n29042 , n6520 , n21665 );
    not g11703 ( n30135 , n12181 );
    xnor g11704 ( n31169 , n7119 , n11272 );
    or g11705 ( n13127 , n14376 , n23051 );
    and g11706 ( n4351 , n23302 , n8663 );
    and g11707 ( n23587 , n11832 , n7616 );
    or g11708 ( n15985 , n11299 , n25286 );
    xnor g11709 ( n22801 , n9971 , n30651 );
    not g11710 ( n2564 , n27031 );
    not g11711 ( n26374 , n14489 );
    not g11712 ( n24387 , n21570 );
    or g11713 ( n716 , n20262 , n14106 );
    and g11714 ( n15595 , n29970 , n30917 );
    xnor g11715 ( n3418 , n4745 , n21137 );
    or g11716 ( n24984 , n24517 , n27789 );
    xnor g11717 ( n13836 , n7289 , n18773 );
    and g11718 ( n12525 , n2468 , n25322 );
    not g11719 ( n16244 , n19317 );
    and g11720 ( n27691 , n3970 , n8594 );
    xnor g11721 ( n19811 , n1141 , n19291 );
    xnor g11722 ( n8083 , n3794 , n3605 );
    xnor g11723 ( n22878 , n21727 , n25386 );
    or g11724 ( n25583 , n5243 , n5248 );
    or g11725 ( n9851 , n30505 , n579 );
    not g11726 ( n30916 , n16077 );
    not g11727 ( n2618 , n891 );
    xor g11728 ( n6182 , n4589 , n1791 );
    or g11729 ( n8554 , n193 , n25738 );
    not g11730 ( n31897 , n16347 );
    and g11731 ( n28883 , n23797 , n710 );
    not g11732 ( n944 , n14954 );
    or g11733 ( n10339 , n6058 , n7307 );
    not g11734 ( n5258 , n15448 );
    or g11735 ( n29931 , n14260 , n23283 );
    nor g11736 ( n14319 , n5022 , n19221 );
    xnor g11737 ( n2540 , n20734 , n14910 );
    nor g11738 ( n13204 , n2001 , n8580 );
    not g11739 ( n19716 , n25444 );
    not g11740 ( n5477 , n9976 );
    and g11741 ( n12258 , n5896 , n5862 );
    xnor g11742 ( n10971 , n29359 , n3567 );
    not g11743 ( n28035 , n15017 );
    and g11744 ( n23878 , n27808 , n28833 );
    xor g11745 ( n18945 , n22779 , n28618 );
    and g11746 ( n7703 , n6411 , n12402 );
    or g11747 ( n9828 , n28332 , n13094 );
    not g11748 ( n1252 , n6972 );
    or g11749 ( n18471 , n14537 , n22345 );
    or g11750 ( n7334 , n1175 , n30253 );
    xor g11751 ( n24777 , n26119 , n6701 );
    not g11752 ( n8152 , n26388 );
    nor g11753 ( n19522 , n7215 , n8172 );
    or g11754 ( n6518 , n4447 , n261 );
    xnor g11755 ( n5295 , n18888 , n4881 );
    not g11756 ( n9282 , n11301 );
    and g11757 ( n8926 , n20617 , n24079 );
    and g11758 ( n22212 , n10907 , n29590 );
    xnor g11759 ( n2264 , n7561 , n9484 );
    xnor g11760 ( n26695 , n7060 , n28277 );
    buf g11761 ( n24601 , n7082 );
    nor g11762 ( n22973 , n3076 , n26639 );
    not g11763 ( n31502 , n21286 );
    xnor g11764 ( n30958 , n2442 , n2075 );
    or g11765 ( n19804 , n18582 , n7223 );
    not g11766 ( n25507 , n2875 );
    xnor g11767 ( n21735 , n6017 , n2632 );
    not g11768 ( n2199 , n10038 );
    xnor g11769 ( n12845 , n25744 , n18817 );
    nor g11770 ( n30980 , n2620 , n14761 );
    xnor g11771 ( n24787 , n7733 , n29697 );
    nor g11772 ( n29111 , n4670 , n13462 );
    xnor g11773 ( n16084 , n8040 , n30158 );
    not g11774 ( n5781 , n5118 );
    nor g11775 ( n30264 , n15153 , n7741 );
    nor g11776 ( n2871 , n26537 , n30369 );
    and g11777 ( n31141 , n7972 , n6841 );
    xnor g11778 ( n9565 , n25593 , n5329 );
    xnor g11779 ( n28303 , n27448 , n14378 );
    xnor g11780 ( n1491 , n4171 , n4407 );
    or g11781 ( n3016 , n8155 , n16269 );
    xnor g11782 ( n26008 , n203 , n3428 );
    xnor g11783 ( n10872 , n5220 , n10474 );
    or g11784 ( n27351 , n26755 , n17960 );
    or g11785 ( n5398 , n23637 , n20361 );
    or g11786 ( n1494 , n29676 , n25988 );
    not g11787 ( n28120 , n3564 );
    not g11788 ( n56 , n18475 );
    not g11789 ( n13247 , n23246 );
    or g11790 ( n15297 , n23607 , n1820 );
    or g11791 ( n23953 , n26663 , n12416 );
    not g11792 ( n13473 , n27201 );
    and g11793 ( n19034 , n19942 , n10114 );
    xor g11794 ( n5267 , n6748 , n7962 );
    not g11795 ( n18080 , n31503 );
    not g11796 ( n17246 , n19345 );
    nor g11797 ( n27234 , n17427 , n24571 );
    and g11798 ( n4245 , n5150 , n445 );
    not g11799 ( n21489 , n6207 );
    and g11800 ( n22176 , n19525 , n30596 );
    xnor g11801 ( n27160 , n23539 , n23381 );
    not g11802 ( n19161 , n20130 );
    or g11803 ( n13692 , n19482 , n14399 );
    and g11804 ( n15825 , n10786 , n6527 );
    or g11805 ( n22340 , n9744 , n29638 );
    xnor g11806 ( n3949 , n602 , n1455 );
    or g11807 ( n2484 , n2231 , n12340 );
    xor g11808 ( n28913 , n18580 , n16283 );
    not g11809 ( n24102 , n19460 );
    and g11810 ( n15968 , n14757 , n20198 );
    xnor g11811 ( n2192 , n13473 , n30949 );
    xnor g11812 ( n29490 , n30795 , n15390 );
    or g11813 ( n29062 , n15288 , n26006 );
    not g11814 ( n5935 , n20359 );
    xnor g11815 ( n21334 , n18253 , n6803 );
    xnor g11816 ( n988 , n7595 , n16437 );
    or g11817 ( n30938 , n3093 , n29776 );
    or g11818 ( n12964 , n3451 , n17372 );
    not g11819 ( n4786 , n11649 );
    and g11820 ( n11511 , n29154 , n22152 );
    and g11821 ( n12051 , n8178 , n12349 );
    not g11822 ( n27918 , n20596 );
    and g11823 ( n5264 , n21938 , n29732 );
    or g11824 ( n14041 , n16841 , n14731 );
    or g11825 ( n1235 , n19615 , n17204 );
    or g11826 ( n10442 , n2395 , n23735 );
    xor g11827 ( n13394 , n25441 , n2070 );
    buf g11828 ( n3570 , n5255 );
    or g11829 ( n30041 , n8561 , n3696 );
    not g11830 ( n23131 , n10463 );
    and g11831 ( n31005 , n8752 , n19380 );
    nor g11832 ( n3767 , n12527 , n8672 );
    or g11833 ( n10906 , n20535 , n19159 );
    not g11834 ( n24620 , n9311 );
    xnor g11835 ( n2603 , n14575 , n15043 );
    or g11836 ( n15084 , n23769 , n17165 );
    nor g11837 ( n19150 , n26429 , n19631 );
    xnor g11838 ( n23455 , n28265 , n10375 );
    xnor g11839 ( n3817 , n4173 , n24479 );
    and g11840 ( n5514 , n23918 , n30060 );
    and g11841 ( n22261 , n1996 , n31118 );
    or g11842 ( n25694 , n248 , n20498 );
    nor g11843 ( n15146 , n25760 , n9239 );
    xnor g11844 ( n4166 , n3616 , n31464 );
    not g11845 ( n27321 , n14691 );
    or g11846 ( n18546 , n8286 , n25412 );
    xnor g11847 ( n1909 , n29213 , n12570 );
    not g11848 ( n6195 , n26996 );
    and g11849 ( n18271 , n1889 , n5150 );
    and g11850 ( n29491 , n20432 , n16735 );
    not g11851 ( n2669 , n26696 );
    xnor g11852 ( n8623 , n4636 , n8217 );
    or g11853 ( n29233 , n27372 , n28539 );
    or g11854 ( n16035 , n29911 , n14428 );
    or g11855 ( n5797 , n30908 , n1375 );
    and g11856 ( n13907 , n16062 , n28176 );
    and g11857 ( n5036 , n15095 , n7098 );
    nor g11858 ( n16866 , n25291 , n19564 );
    not g11859 ( n1022 , n13648 );
    not g11860 ( n399 , n4828 );
    or g11861 ( n18111 , n18584 , n6547 );
    not g11862 ( n23983 , n13488 );
    xnor g11863 ( n31254 , n5617 , n6066 );
    not g11864 ( n26773 , n11660 );
    or g11865 ( n25836 , n2862 , n3604 );
    not g11866 ( n3595 , n24833 );
    not g11867 ( n12621 , n9835 );
    not g11868 ( n20558 , n4586 );
    or g11869 ( n11276 , n27348 , n15074 );
    and g11870 ( n12292 , n11077 , n17167 );
    not g11871 ( n28527 , n13454 );
    not g11872 ( n17426 , n3979 );
    nor g11873 ( n20997 , n3837 , n14925 );
    and g11874 ( n27394 , n12722 , n254 );
    or g11875 ( n644 , n27883 , n14136 );
    or g11876 ( n3518 , n4067 , n20233 );
    not g11877 ( n17960 , n16054 );
    or g11878 ( n28702 , n15444 , n3187 );
    not g11879 ( n24710 , n14842 );
    not g11880 ( n25771 , n11561 );
    or g11881 ( n31180 , n14020 , n1790 );
    or g11882 ( n15486 , n24988 , n6800 );
    not g11883 ( n25259 , n2170 );
    xnor g11884 ( n29705 , n8463 , n14466 );
    and g11885 ( n373 , n7866 , n5374 );
    or g11886 ( n5259 , n1803 , n17998 );
    or g11887 ( n2499 , n27087 , n23708 );
    and g11888 ( n23854 , n30770 , n31399 );
    and g11889 ( n10665 , n24254 , n2678 );
    not g11890 ( n13346 , n28158 );
    or g11891 ( n6059 , n5469 , n9432 );
    not g11892 ( n25399 , n5075 );
    not g11893 ( n7729 , n974 );
    xnor g11894 ( n27284 , n21388 , n18839 );
    or g11895 ( n18320 , n28806 , n6210 );
    or g11896 ( n1826 , n16367 , n30094 );
    not g11897 ( n3509 , n10034 );
    xnor g11898 ( n14599 , n7380 , n17376 );
    and g11899 ( n23940 , n11657 , n10080 );
    not g11900 ( n2372 , n24361 );
    not g11901 ( n12446 , n23628 );
    or g11902 ( n18556 , n8489 , n17087 );
    or g11903 ( n27519 , n4931 , n25307 );
    or g11904 ( n3608 , n5422 , n17223 );
    not g11905 ( n5410 , n17100 );
    or g11906 ( n27198 , n24699 , n24285 );
    xnor g11907 ( n25378 , n30851 , n20522 );
    not g11908 ( n15125 , n18866 );
    or g11909 ( n8903 , n28479 , n27675 );
    xnor g11910 ( n6986 , n14226 , n25214 );
    and g11911 ( n17276 , n9817 , n6514 );
    xnor g11912 ( n7557 , n26210 , n30096 );
    xnor g11913 ( n5860 , n7897 , n3996 );
    not g11914 ( n24643 , n15854 );
    not g11915 ( n23263 , n9061 );
    xnor g11916 ( n16079 , n31760 , n3783 );
    not g11917 ( n21066 , n7999 );
    not g11918 ( n2513 , n13992 );
    and g11919 ( n23721 , n14433 , n6677 );
    not g11920 ( n2007 , n26630 );
    xor g11921 ( n5055 , n21281 , n26033 );
    or g11922 ( n30857 , n18232 , n15973 );
    or g11923 ( n13673 , n7367 , n17678 );
    xnor g11924 ( n30246 , n4588 , n25724 );
    nor g11925 ( n16621 , n9116 , n30934 );
    xnor g11926 ( n14195 , n2572 , n4276 );
    not g11927 ( n12222 , n13221 );
    not g11928 ( n21869 , n21778 );
    and g11929 ( n19813 , n30592 , n21294 );
    and g11930 ( n19657 , n30417 , n7036 );
    and g11931 ( n446 , n12357 , n19689 );
    not g11932 ( n12762 , n7728 );
    xnor g11933 ( n29990 , n22795 , n22148 );
    not g11934 ( n20996 , n21089 );
    not g11935 ( n19134 , n16384 );
    not g11936 ( n1396 , n5616 );
    xnor g11937 ( n25555 , n20014 , n18439 );
    xnor g11938 ( n2242 , n21610 , n1366 );
    and g11939 ( n10985 , n28473 , n16009 );
    not g11940 ( n3738 , n11791 );
    not g11941 ( n24518 , n2558 );
    buf g11942 ( n22248 , n12178 );
    not g11943 ( n10601 , n318 );
    xnor g11944 ( n27524 , n14619 , n6604 );
    or g11945 ( n19323 , n12654 , n12458 );
    or g11946 ( n6011 , n23891 , n2190 );
    xnor g11947 ( n6040 , n10618 , n4026 );
    not g11948 ( n18164 , n30921 );
    not g11949 ( n10090 , n18177 );
    not g11950 ( n26328 , n21263 );
    not g11951 ( n14132 , n26632 );
    not g11952 ( n26956 , n4106 );
    and g11953 ( n5426 , n7309 , n13273 );
    nor g11954 ( n1086 , n10338 , n12318 );
    not g11955 ( n2106 , n18837 );
    xnor g11956 ( n31784 , n11156 , n21412 );
    and g11957 ( n24328 , n20925 , n1514 );
    not g11958 ( n4424 , n23839 );
    xnor g11959 ( n19260 , n19632 , n24137 );
    not g11960 ( n20369 , n1689 );
    not g11961 ( n8747 , n21979 );
    or g11962 ( n2789 , n15384 , n16965 );
    xor g11963 ( n5108 , n4691 , n10612 );
    xnor g11964 ( n16807 , n19733 , n3793 );
    and g11965 ( n15800 , n24949 , n22226 );
    or g11966 ( n7935 , n17212 , n15781 );
    or g11967 ( n27926 , n20157 , n20744 );
    and g11968 ( n31858 , n26450 , n11326 );
    xnor g11969 ( n24826 , n18736 , n11209 );
    xnor g11970 ( n12653 , n1919 , n11076 );
    or g11971 ( n24342 , n10460 , n21668 );
    xnor g11972 ( n23789 , n16330 , n9088 );
    not g11973 ( n22804 , n5989 );
    and g11974 ( n16371 , n24284 , n19723 );
    or g11975 ( n349 , n28935 , n20777 );
    and g11976 ( n28051 , n490 , n9581 );
    xnor g11977 ( n19901 , n8561 , n24578 );
    xnor g11978 ( n5125 , n31363 , n175 );
    not g11979 ( n27919 , n19255 );
    not g11980 ( n13503 , n23983 );
    or g11981 ( n15184 , n23889 , n23187 );
    and g11982 ( n14126 , n23227 , n14032 );
    xor g11983 ( n11725 , n7110 , n8201 );
    nor g11984 ( n1873 , n17166 , n24401 );
    or g11985 ( n6865 , n5300 , n3484 );
    xnor g11986 ( n20904 , n18583 , n28914 );
    nor g11987 ( n18741 , n24003 , n17985 );
    or g11988 ( n7266 , n24704 , n22019 );
    not g11989 ( n31894 , n14612 );
    and g11990 ( n18463 , n20508 , n29910 );
    and g11991 ( n2442 , n6802 , n30755 );
    nor g11992 ( n13770 , n1995 , n12319 );
    or g11993 ( n21990 , n8804 , n27716 );
    or g11994 ( n6237 , n21136 , n27715 );
    xnor g11995 ( n21816 , n22157 , n21466 );
    not g11996 ( n19916 , n13971 );
    xnor g11997 ( n29265 , n31550 , n26301 );
    not g11998 ( n5905 , n11935 );
    nor g11999 ( n11075 , n20799 , n3039 );
    xnor g12000 ( n27364 , n21330 , n3850 );
    or g12001 ( n26513 , n11385 , n23820 );
    not g12002 ( n27457 , n15828 );
    not g12003 ( n15568 , n7434 );
    or g12004 ( n4094 , n19431 , n19912 );
    buf g12005 ( n9486 , n30174 );
    or g12006 ( n9405 , n5400 , n11760 );
    not g12007 ( n15593 , n22855 );
    xnor g12008 ( n10288 , n27673 , n1965 );
    xnor g12009 ( n869 , n26995 , n18417 );
    or g12010 ( n4359 , n10393 , n28026 );
    or g12011 ( n25611 , n17484 , n24545 );
    not g12012 ( n2512 , n19902 );
    not g12013 ( n13159 , n10367 );
    not g12014 ( n831 , n4606 );
    xnor g12015 ( n3257 , n13553 , n8052 );
    nor g12016 ( n28487 , n9963 , n27167 );
    xnor g12017 ( n31787 , n25923 , n1274 );
    and g12018 ( n28515 , n11933 , n320 );
    and g12019 ( n10309 , n7282 , n14197 );
    and g12020 ( n7681 , n15553 , n20792 );
    or g12021 ( n16699 , n7654 , n5353 );
    xnor g12022 ( n8462 , n4250 , n1966 );
    or g12023 ( n23436 , n13631 , n21437 );
    or g12024 ( n20458 , n52 , n13747 );
    or g12025 ( n17139 , n4508 , n3749 );
    xnor g12026 ( n13710 , n11529 , n1272 );
    not g12027 ( n4458 , n25358 );
    and g12028 ( n10822 , n31795 , n13362 );
    or g12029 ( n578 , n4664 , n12094 );
    not g12030 ( n13101 , n10860 );
    or g12031 ( n18797 , n19427 , n10108 );
    xnor g12032 ( n6066 , n20769 , n3030 );
    nor g12033 ( n22186 , n15864 , n3258 );
    not g12034 ( n2712 , n7314 );
    nor g12035 ( n22947 , n20262 , n26961 );
    xnor g12036 ( n17376 , n30560 , n22092 );
    or g12037 ( n15171 , n23764 , n16234 );
    or g12038 ( n7462 , n28364 , n11277 );
    or g12039 ( n1651 , n23884 , n19845 );
    xnor g12040 ( n22371 , n17372 , n11293 );
    not g12041 ( n13945 , n5108 );
    xnor g12042 ( n15805 , n9064 , n24008 );
    not g12043 ( n14194 , n19283 );
    xnor g12044 ( n17527 , n27878 , n9122 );
    not g12045 ( n6685 , n26616 );
    or g12046 ( n26730 , n25950 , n26337 );
    not g12047 ( n20517 , n15357 );
    xnor g12048 ( n946 , n12937 , n3186 );
    not g12049 ( n4443 , n4627 );
    or g12050 ( n7306 , n30875 , n16915 );
    or g12051 ( n21734 , n15595 , n17637 );
    xnor g12052 ( n27271 , n23175 , n15901 );
    not g12053 ( n3706 , n29933 );
    or g12054 ( n9112 , n14455 , n31478 );
    or g12055 ( n16372 , n22724 , n27099 );
    not g12056 ( n1343 , n28458 );
    and g12057 ( n12081 , n26175 , n20919 );
    and g12058 ( n31997 , n14863 , n22949 );
    not g12059 ( n7541 , n20109 );
    nor g12060 ( n15719 , n28394 , n31773 );
    xnor g12061 ( n16933 , n15696 , n23357 );
    not g12062 ( n5419 , n8536 );
    xnor g12063 ( n4650 , n24972 , n17901 );
    or g12064 ( n24292 , n15816 , n17809 );
    not g12065 ( n7087 , n29484 );
    or g12066 ( n17397 , n24163 , n13625 );
    xnor g12067 ( n8058 , n6731 , n5895 );
    buf g12068 ( n23735 , n24676 );
    or g12069 ( n2661 , n9891 , n406 );
    xnor g12070 ( n30296 , n12119 , n30067 );
    nor g12071 ( n1756 , n13210 , n20644 );
    and g12072 ( n8789 , n15481 , n27934 );
    and g12073 ( n20552 , n26554 , n7266 );
    xnor g12074 ( n4433 , n1179 , n10875 );
    and g12075 ( n25082 , n23712 , n14698 );
    not g12076 ( n10444 , n10040 );
    or g12077 ( n23950 , n30326 , n27534 );
    and g12078 ( n9498 , n2544 , n7241 );
    and g12079 ( n2171 , n10104 , n30287 );
    or g12080 ( n28657 , n12882 , n27695 );
    nor g12081 ( n6335 , n20862 , n3030 );
    or g12082 ( n10173 , n14264 , n7515 );
    or g12083 ( n22116 , n19973 , n453 );
    not g12084 ( n1957 , n19105 );
    xnor g12085 ( n29640 , n12938 , n31426 );
    or g12086 ( n2391 , n31720 , n22680 );
    xnor g12087 ( n7193 , n8396 , n19775 );
    xnor g12088 ( n15012 , n3837 , n14925 );
    and g12089 ( n19001 , n13782 , n2740 );
    or g12090 ( n11122 , n3357 , n16433 );
    not g12091 ( n29810 , n21716 );
    xnor g12092 ( n23409 , n15276 , n20695 );
    nor g12093 ( n3529 , n29946 , n28940 );
    xnor g12094 ( n20475 , n5707 , n1584 );
    and g12095 ( n27424 , n659 , n1884 );
    not g12096 ( n3110 , n9801 );
    xnor g12097 ( n29102 , n9039 , n11729 );
    xnor g12098 ( n13723 , n29358 , n5014 );
    nor g12099 ( n31029 , n28305 , n350 );
    and g12100 ( n29813 , n2107 , n667 );
    not g12101 ( n29982 , n15750 );
    or g12102 ( n8218 , n2219 , n5763 );
    not g12103 ( n8558 , n11306 );
    nor g12104 ( n24474 , n31783 , n21508 );
    xor g12105 ( n4048 , n14614 , n1320 );
    or g12106 ( n14550 , n17876 , n4366 );
    xnor g12107 ( n29763 , n1959 , n17501 );
    xnor g12108 ( n18167 , n11360 , n17109 );
    not g12109 ( n27176 , n1529 );
    not g12110 ( n10837 , n18842 );
    not g12111 ( n30218 , n14410 );
    not g12112 ( n13515 , n21168 );
    and g12113 ( n17707 , n9767 , n23894 );
    not g12114 ( n16683 , n28242 );
    or g12115 ( n5214 , n10029 , n8018 );
    and g12116 ( n9264 , n8799 , n16348 );
    nor g12117 ( n14056 , n29764 , n14696 );
    xnor g12118 ( n25156 , n26894 , n22867 );
    or g12119 ( n2281 , n15085 , n25503 );
    xnor g12120 ( n10884 , n11373 , n19405 );
    xnor g12121 ( n19312 , n29419 , n25058 );
    not g12122 ( n3403 , n7655 );
    xnor g12123 ( n16651 , n10667 , n6517 );
    xnor g12124 ( n6792 , n2612 , n9772 );
    xnor g12125 ( n2173 , n30965 , n20034 );
    xnor g12126 ( n3585 , n26991 , n31338 );
    not g12127 ( n16 , n10244 );
    xnor g12128 ( n8381 , n28267 , n10451 );
    not g12129 ( n19350 , n28325 );
    not g12130 ( n7122 , n19622 );
    xnor g12131 ( n7310 , n22279 , n26786 );
    nor g12132 ( n24048 , n10423 , n2808 );
    and g12133 ( n26444 , n31304 , n28657 );
    not g12134 ( n26977 , n14795 );
    and g12135 ( n6941 , n27189 , n9295 );
    or g12136 ( n11784 , n9072 , n8818 );
    not g12137 ( n16399 , n4201 );
    and g12138 ( n19616 , n27597 , n11927 );
    not g12139 ( n27101 , n14825 );
    xnor g12140 ( n30150 , n14186 , n27422 );
    xor g12141 ( n8579 , n29012 , n21906 );
    and g12142 ( n10212 , n26850 , n19284 );
    xnor g12143 ( n20386 , n3592 , n1856 );
    not g12144 ( n21023 , n7872 );
    not g12145 ( n25154 , n11250 );
    xnor g12146 ( n17675 , n29146 , n17387 );
    nor g12147 ( n7120 , n20151 , n23004 );
    not g12148 ( n14123 , n13259 );
    not g12149 ( n31 , n23994 );
    xnor g12150 ( n7844 , n17546 , n2629 );
    not g12151 ( n21513 , n10338 );
    xnor g12152 ( n30064 , n26723 , n21768 );
    not g12153 ( n26623 , n2014 );
    xnor g12154 ( n27713 , n13856 , n26573 );
    xnor g12155 ( n1694 , n5388 , n18002 );
    not g12156 ( n28976 , n31884 );
    or g12157 ( n3819 , n22158 , n22953 );
    or g12158 ( n4251 , n30618 , n16355 );
    nor g12159 ( n95 , n5441 , n21390 );
    and g12160 ( n28982 , n29757 , n5000 );
    nor g12161 ( n99 , n4093 , n4012 );
    xnor g12162 ( n21642 , n21248 , n12955 );
    xnor g12163 ( n23663 , n23184 , n26203 );
    or g12164 ( n9606 , n25801 , n27084 );
    or g12165 ( n9995 , n18545 , n29374 );
    and g12166 ( n8178 , n29964 , n28089 );
    not g12167 ( n28002 , n11903 );
    or g12168 ( n31796 , n27527 , n29280 );
    xnor g12169 ( n11992 , n27034 , n26758 );
    and g12170 ( n16355 , n18642 , n1542 );
    not g12171 ( n894 , n24691 );
    not g12172 ( n4765 , n30541 );
    xnor g12173 ( n27935 , n21159 , n19619 );
    nor g12174 ( n30701 , n20588 , n30812 );
    or g12175 ( n17258 , n12309 , n11391 );
    or g12176 ( n27964 , n20983 , n2440 );
    xnor g12177 ( n634 , n23195 , n30287 );
    xnor g12178 ( n4947 , n9662 , n18236 );
    xnor g12179 ( n31836 , n24921 , n8747 );
    and g12180 ( n17742 , n15889 , n1499 );
    or g12181 ( n24339 , n24426 , n18898 );
    not g12182 ( n14533 , n231 );
    nor g12183 ( n25408 , n29039 , n19002 );
    not g12184 ( n15288 , n29249 );
    nor g12185 ( n31454 , n12237 , n27811 );
    and g12186 ( n15969 , n12846 , n681 );
    and g12187 ( n9700 , n12452 , n11020 );
    and g12188 ( n10667 , n23808 , n9030 );
    not g12189 ( n24624 , n4767 );
    not g12190 ( n21314 , n6349 );
    and g12191 ( n18437 , n7067 , n5424 );
    nor g12192 ( n20143 , n8518 , n14768 );
    xnor g12193 ( n3370 , n30305 , n23511 );
    not g12194 ( n29245 , n12222 );
    or g12195 ( n15230 , n23770 , n20533 );
    or g12196 ( n16632 , n22711 , n14304 );
    or g12197 ( n31385 , n17696 , n24835 );
    xnor g12198 ( n17720 , n6445 , n17913 );
    not g12199 ( n15795 , n2334 );
    buf g12200 ( n14558 , n5706 );
    not g12201 ( n28360 , n18751 );
    not g12202 ( n15346 , n2741 );
    xnor g12203 ( n27187 , n28410 , n31060 );
    not g12204 ( n5709 , n19256 );
    or g12205 ( n12736 , n25366 , n16314 );
    xnor g12206 ( n6424 , n16627 , n7830 );
    not g12207 ( n23991 , n2199 );
    and g12208 ( n24843 , n26081 , n31656 );
    not g12209 ( n227 , n21342 );
    and g12210 ( n12071 , n31699 , n9314 );
    xnor g12211 ( n18424 , n31667 , n31887 );
    or g12212 ( n31666 , n10034 , n17898 );
    and g12213 ( n19490 , n1844 , n19959 );
    xnor g12214 ( n5057 , n29324 , n26496 );
    xnor g12215 ( n29006 , n3907 , n15749 );
    xnor g12216 ( n5379 , n20642 , n19524 );
    xnor g12217 ( n15320 , n23278 , n3259 );
    xor g12218 ( n26694 , n23022 , n24649 );
    xnor g12219 ( n30259 , n21860 , n12972 );
    xnor g12220 ( n20800 , n19181 , n1353 );
    xnor g12221 ( n15807 , n18226 , n4977 );
    or g12222 ( n422 , n20413 , n25612 );
    not g12223 ( n31067 , n13831 );
    xnor g12224 ( n27716 , n3638 , n3289 );
    and g12225 ( n14325 , n19157 , n19172 );
    xnor g12226 ( n19044 , n15217 , n31339 );
    not g12227 ( n28566 , n15159 );
    not g12228 ( n25159 , n766 );
    and g12229 ( n13732 , n19874 , n16508 );
    not g12230 ( n28357 , n17638 );
    nor g12231 ( n23576 , n28559 , n12899 );
    or g12232 ( n786 , n17362 , n30891 );
    not g12233 ( n27143 , n25843 );
    or g12234 ( n5713 , n29257 , n14314 );
    and g12235 ( n11164 , n14991 , n168 );
    xnor g12236 ( n21703 , n14248 , n5452 );
    and g12237 ( n10472 , n22617 , n11464 );
    not g12238 ( n190 , n4907 );
    nor g12239 ( n21400 , n28978 , n11716 );
    not g12240 ( n5165 , n6564 );
    or g12241 ( n31779 , n10539 , n15478 );
    not g12242 ( n12349 , n17068 );
    not g12243 ( n1232 , n397 );
    and g12244 ( n5019 , n8056 , n17766 );
    nor g12245 ( n16039 , n4918 , n11815 );
    not g12246 ( n10532 , n14004 );
    nor g12247 ( n17423 , n16157 , n22126 );
    and g12248 ( n7652 , n10903 , n716 );
    xnor g12249 ( n24669 , n9199 , n26656 );
    xnor g12250 ( n12672 , n31420 , n22580 );
    xnor g12251 ( n17039 , n5435 , n1331 );
    xnor g12252 ( n6470 , n5990 , n14044 );
    xnor g12253 ( n27320 , n2346 , n6826 );
    not g12254 ( n15792 , n13332 );
    xnor g12255 ( n28890 , n11594 , n31595 );
    nor g12256 ( n968 , n30434 , n12108 );
    not g12257 ( n13067 , n31310 );
    and g12258 ( n30324 , n25905 , n19884 );
    or g12259 ( n16507 , n23358 , n16452 );
    and g12260 ( n17799 , n1512 , n11117 );
    xnor g12261 ( n28636 , n13511 , n27320 );
    nor g12262 ( n19514 , n16836 , n14844 );
    not g12263 ( n25728 , n30425 );
    xnor g12264 ( n14076 , n22542 , n17099 );
    not g12265 ( n23096 , n3086 );
    and g12266 ( n19469 , n19483 , n9236 );
    xnor g12267 ( n7508 , n4832 , n6707 );
    and g12268 ( n17067 , n15243 , n1428 );
    xnor g12269 ( n4412 , n10983 , n10610 );
    and g12270 ( n3833 , n2633 , n31385 );
    not g12271 ( n4427 , n24464 );
    xnor g12272 ( n24716 , n10008 , n15262 );
    not g12273 ( n5013 , n27360 );
    xnor g12274 ( n1601 , n17617 , n5069 );
    xnor g12275 ( n22107 , n31644 , n19273 );
    not g12276 ( n10058 , n26163 );
    or g12277 ( n28729 , n17971 , n2007 );
    not g12278 ( n3192 , n26137 );
    or g12279 ( n26320 , n5733 , n25579 );
    not g12280 ( n29777 , n1010 );
    xnor g12281 ( n7730 , n18349 , n2693 );
    or g12282 ( n20461 , n16200 , n73 );
    or g12283 ( n32013 , n19255 , n29400 );
    not g12284 ( n29851 , n10395 );
    not g12285 ( n27763 , n25793 );
    and g12286 ( n5630 , n18636 , n19964 );
    xnor g12287 ( n20308 , n20654 , n3633 );
    or g12288 ( n11809 , n2044 , n25587 );
    not g12289 ( n21547 , n24414 );
    or g12290 ( n11459 , n14951 , n756 );
    not g12291 ( n6910 , n18518 );
    not g12292 ( n8975 , n31424 );
    or g12293 ( n18716 , n15329 , n11525 );
    not g12294 ( n17642 , n24995 );
    not g12295 ( n9395 , n28998 );
    and g12296 ( n28698 , n7221 , n16554 );
    and g12297 ( n28844 , n12014 , n7473 );
    not g12298 ( n8555 , n1730 );
    not g12299 ( n30003 , n23633 );
    not g12300 ( n13405 , n8600 );
    xnor g12301 ( n27962 , n9321 , n25805 );
    not g12302 ( n20796 , n12412 );
    or g12303 ( n29312 , n1371 , n2409 );
    and g12304 ( n5619 , n25923 , n6237 );
    not g12305 ( n15778 , n2408 );
    not g12306 ( n8601 , n10073 );
    xnor g12307 ( n9727 , n24132 , n23400 );
    or g12308 ( n18178 , n26705 , n26006 );
    or g12309 ( n26167 , n17255 , n14437 );
    or g12310 ( n15350 , n25800 , n10526 );
    and g12311 ( n11342 , n2426 , n22284 );
    xnor g12312 ( n9592 , n20262 , n14106 );
    not g12313 ( n10893 , n8910 );
    xnor g12314 ( n5546 , n18551 , n12777 );
    and g12315 ( n19448 , n3732 , n14793 );
    not g12316 ( n13729 , n6819 );
    and g12317 ( n21952 , n28711 , n27942 );
    or g12318 ( n10586 , n3203 , n4745 );
    or g12319 ( n2584 , n4264 , n24121 );
    xnor g12320 ( n22865 , n18720 , n2095 );
    xnor g12321 ( n31888 , n10773 , n20236 );
    or g12322 ( n21611 , n19138 , n29367 );
    not g12323 ( n12841 , n11747 );
    nor g12324 ( n2286 , n20017 , n11913 );
    not g12325 ( n24343 , n7014 );
    or g12326 ( n9903 , n23784 , n3251 );
    not g12327 ( n14134 , n19056 );
    xnor g12328 ( n24800 , n16292 , n2610 );
    not g12329 ( n4890 , n12388 );
    not g12330 ( n27906 , n12998 );
    not g12331 ( n10050 , n11921 );
    and g12332 ( n5239 , n23242 , n25622 );
    not g12333 ( n673 , n31258 );
    and g12334 ( n27425 , n17838 , n19473 );
    xnor g12335 ( n3475 , n25067 , n4631 );
    xnor g12336 ( n6250 , n10009 , n22827 );
    and g12337 ( n649 , n896 , n8935 );
    nor g12338 ( n8302 , n7180 , n24578 );
    not g12339 ( n18191 , n21928 );
    not g12340 ( n17142 , n30887 );
    or g12341 ( n17202 , n14276 , n18670 );
    xnor g12342 ( n477 , n25525 , n3407 );
    xnor g12343 ( n19371 , n4852 , n12223 );
    not g12344 ( n18902 , n3029 );
    not g12345 ( n8585 , n31940 );
    xnor g12346 ( n14839 , n13217 , n22679 );
    xnor g12347 ( n6810 , n18384 , n27534 );
    and g12348 ( n30583 , n24543 , n1135 );
    and g12349 ( n17483 , n17659 , n13078 );
    and g12350 ( n29835 , n29758 , n24799 );
    and g12351 ( n9201 , n19895 , n10935 );
    not g12352 ( n7767 , n20135 );
    and g12353 ( n3723 , n16336 , n26310 );
    not g12354 ( n18257 , n31711 );
    nor g12355 ( n13883 , n23061 , n2169 );
    and g12356 ( n23102 , n13442 , n2670 );
    not g12357 ( n4202 , n10904 );
    and g12358 ( n438 , n16460 , n11848 );
    not g12359 ( n21768 , n10084 );
    not g12360 ( n29422 , n17382 );
    or g12361 ( n8185 , n5447 , n905 );
    xnor g12362 ( n4848 , n21936 , n21459 );
    xnor g12363 ( n5241 , n19034 , n3527 );
    and g12364 ( n22080 , n11081 , n22674 );
    xnor g12365 ( n8239 , n12739 , n12399 );
    xnor g12366 ( n13667 , n6420 , n6778 );
    or g12367 ( n23711 , n1177 , n25130 );
    and g12368 ( n24705 , n8060 , n9142 );
    not g12369 ( n19983 , n27743 );
    nor g12370 ( n25879 , n20495 , n6331 );
    not g12371 ( n9612 , n15593 );
    or g12372 ( n31574 , n6534 , n4525 );
    xnor g12373 ( n27630 , n16882 , n22361 );
    not g12374 ( n24908 , n18652 );
    xnor g12375 ( n13683 , n5948 , n20390 );
    or g12376 ( n8055 , n25282 , n24602 );
    not g12377 ( n58 , n24360 );
    not g12378 ( n12582 , n8013 );
    xnor g12379 ( n10696 , n3560 , n16401 );
    and g12380 ( n27142 , n8942 , n8825 );
    and g12381 ( n5682 , n7384 , n14902 );
    xnor g12382 ( n8666 , n28075 , n14338 );
    or g12383 ( n8957 , n7895 , n10648 );
    nor g12384 ( n27655 , n7465 , n6819 );
    and g12385 ( n2702 , n25056 , n3863 );
    and g12386 ( n7289 , n24986 , n23420 );
    xnor g12387 ( n29173 , n22928 , n16786 );
    not g12388 ( n28884 , n7588 );
    xnor g12389 ( n29141 , n21828 , n13683 );
    not g12390 ( n31988 , n16462 );
    not g12391 ( n5779 , n3910 );
    xnor g12392 ( n8335 , n9116 , n18388 );
    or g12393 ( n21479 , n3529 , n5318 );
    or g12394 ( n13891 , n20352 , n18646 );
    xnor g12395 ( n26153 , n21215 , n23605 );
    and g12396 ( n19821 , n19521 , n21673 );
    not g12397 ( n16979 , n21244 );
    or g12398 ( n2738 , n24745 , n6898 );
    xnor g12399 ( n31570 , n6572 , n15723 );
    xnor g12400 ( n7910 , n20495 , n7209 );
    not g12401 ( n4192 , n21712 );
    not g12402 ( n8704 , n14260 );
    not g12403 ( n208 , n17834 );
    not g12404 ( n1230 , n25169 );
    xnor g12405 ( n2506 , n1935 , n23681 );
    xnor g12406 ( n8369 , n3946 , n27264 );
    not g12407 ( n19922 , n12123 );
    or g12408 ( n7673 , n7014 , n7408 );
    or g12409 ( n957 , n12324 , n29563 );
    and g12410 ( n30621 , n7550 , n20230 );
    xnor g12411 ( n1827 , n15306 , n25702 );
    not g12412 ( n27787 , n1518 );
    or g12413 ( n19826 , n24877 , n1264 );
    or g12414 ( n10850 , n7570 , n3161 );
    not g12415 ( n15450 , n631 );
    xnor g12416 ( n17313 , n13458 , n25848 );
    not g12417 ( n23722 , n22015 );
    and g12418 ( n28737 , n10886 , n6374 );
    not g12419 ( n1381 , n22721 );
    not g12420 ( n24235 , n14385 );
    or g12421 ( n15483 , n21396 , n2634 );
    xnor g12422 ( n12204 , n13454 , n30458 );
    xnor g12423 ( n18710 , n20870 , n26636 );
    and g12424 ( n20348 , n15872 , n14562 );
    xor g12425 ( n25210 , n20068 , n29101 );
    not g12426 ( n6861 , n17454 );
    not g12427 ( n6538 , n2746 );
    not g12428 ( n6552 , n13800 );
    not g12429 ( n18133 , n17986 );
    nor g12430 ( n15529 , n23915 , n2260 );
    or g12431 ( n27759 , n20632 , n20759 );
    or g12432 ( n10745 , n14302 , n10234 );
    nor g12433 ( n31582 , n16312 , n22109 );
    or g12434 ( n18488 , n27123 , n22682 );
    buf g12435 ( n7017 , n10684 );
    nor g12436 ( n26036 , n20510 , n19716 );
    xnor g12437 ( n21945 , n19002 , n8988 );
    and g12438 ( n8034 , n27265 , n12336 );
    not g12439 ( n31259 , n18518 );
    or g12440 ( n98 , n29132 , n22924 );
    xor g12441 ( n3367 , n24232 , n27974 );
    and g12442 ( n3083 , n18906 , n31738 );
    or g12443 ( n14164 , n5130 , n23333 );
    xnor g12444 ( n16927 , n9129 , n29322 );
    or g12445 ( n2517 , n11406 , n31714 );
    not g12446 ( n10622 , n12897 );
    xnor g12447 ( n2521 , n25390 , n29528 );
    and g12448 ( n17155 , n23759 , n13819 );
    nor g12449 ( n688 , n18253 , n22075 );
    or g12450 ( n25664 , n2754 , n30319 );
    and g12451 ( n8887 , n16682 , n23450 );
    not g12452 ( n2023 , n29046 );
    not g12453 ( n10537 , n21956 );
    not g12454 ( n8119 , n31028 );
    not g12455 ( n27956 , n29346 );
    or g12456 ( n22444 , n13530 , n12059 );
    not g12457 ( n14018 , n4021 );
    xnor g12458 ( n6546 , n19677 , n25467 );
    or g12459 ( n686 , n25154 , n13336 );
    xnor g12460 ( n6924 , n2582 , n11949 );
    or g12461 ( n2659 , n2184 , n8669 );
    and g12462 ( n17779 , n16218 , n3254 );
    xnor g12463 ( n16190 , n21597 , n30411 );
    and g12464 ( n16695 , n9425 , n11591 );
    or g12465 ( n28000 , n21408 , n29462 );
    not g12466 ( n26322 , n31873 );
    nor g12467 ( n28191 , n3080 , n22493 );
    nor g12468 ( n13052 , n11065 , n3692 );
    not g12469 ( n24871 , n17918 );
    and g12470 ( n20868 , n21460 , n5236 );
    or g12471 ( n27296 , n3640 , n29900 );
    or g12472 ( n16691 , n30680 , n14169 );
    xnor g12473 ( n16324 , n22805 , n26037 );
    not g12474 ( n7979 , n7541 );
    not g12475 ( n18772 , n22181 );
    nor g12476 ( n15446 , n21197 , n12604 );
    not g12477 ( n12543 , n11049 );
    not g12478 ( n24457 , n20192 );
    xor g12479 ( n20312 , n23664 , n21429 );
    xnor g12480 ( n22178 , n21641 , n18910 );
    or g12481 ( n19091 , n14356 , n6985 );
    xnor g12482 ( n134 , n954 , n12991 );
    or g12483 ( n12791 , n3847 , n102 );
    nor g12484 ( n20671 , n7414 , n26423 );
    and g12485 ( n29618 , n18987 , n26915 );
    nor g12486 ( n18916 , n4350 , n24056 );
    and g12487 ( n4660 , n32022 , n10225 );
    xor g12488 ( n9566 , n11904 , n23198 );
    nor g12489 ( n10691 , n23115 , n28453 );
    xnor g12490 ( n6183 , n10707 , n5948 );
    xnor g12491 ( n26765 , n27575 , n10334 );
    and g12492 ( n27728 , n16398 , n12918 );
    nor g12493 ( n3648 , n27972 , n21735 );
    not g12494 ( n26061 , n11035 );
    not g12495 ( n20140 , n17906 );
    and g12496 ( n6598 , n2738 , n16748 );
    or g12497 ( n21645 , n22002 , n31977 );
    or g12498 ( n17297 , n28467 , n16207 );
    not g12499 ( n3587 , n14134 );
    or g12500 ( n9319 , n19931 , n23155 );
    xnor g12501 ( n1433 , n26930 , n5635 );
    not g12502 ( n18653 , n23183 );
    or g12503 ( n3886 , n20576 , n16349 );
    xnor g12504 ( n25480 , n16304 , n1720 );
    xnor g12505 ( n18620 , n18900 , n6861 );
    or g12506 ( n21101 , n22446 , n30183 );
    nor g12507 ( n20139 , n19494 , n27531 );
    not g12508 ( n8506 , n17149 );
    xnor g12509 ( n24738 , n14339 , n13767 );
    or g12510 ( n7837 , n20231 , n22503 );
    xnor g12511 ( n523 , n16094 , n7843 );
    or g12512 ( n17238 , n20881 , n15589 );
    or g12513 ( n22068 , n1801 , n10596 );
    not g12514 ( n29695 , n3154 );
    not g12515 ( n24733 , n24991 );
    and g12516 ( n13730 , n25744 , n5698 );
    xnor g12517 ( n13540 , n27608 , n30830 );
    nor g12518 ( n18455 , n24191 , n10860 );
    or g12519 ( n24142 , n19838 , n639 );
    not g12520 ( n11341 , n13137 );
    xnor g12521 ( n13837 , n15309 , n24455 );
    nor g12522 ( n24571 , n11723 , n11093 );
    or g12523 ( n12466 , n2957 , n2771 );
    not g12524 ( n18827 , n24537 );
    or g12525 ( n5437 , n28008 , n13527 );
    not g12526 ( n10153 , n30141 );
    or g12527 ( n16627 , n2252 , n4888 );
    and g12528 ( n12457 , n9926 , n19272 );
    xnor g12529 ( n28541 , n27295 , n6087 );
    not g12530 ( n3029 , n15671 );
    xnor g12531 ( n4021 , n30048 , n2545 );
    and g12532 ( n28279 , n15705 , n16464 );
    nor g12533 ( n6092 , n12139 , n6014 );
    or g12534 ( n1083 , n8075 , n15962 );
    and g12535 ( n5891 , n3217 , n27825 );
    not g12536 ( n20431 , n7582 );
    not g12537 ( n11117 , n21392 );
    nor g12538 ( n18247 , n18645 , n23306 );
    not g12539 ( n24362 , n10737 );
    not g12540 ( n4973 , n30964 );
    and g12541 ( n14482 , n4912 , n9158 );
    not g12542 ( n31627 , n19410 );
    or g12543 ( n28861 , n2573 , n7505 );
    or g12544 ( n23193 , n721 , n24266 );
    xnor g12545 ( n23557 , n14819 , n19771 );
    xnor g12546 ( n23582 , n17149 , n20881 );
    or g12547 ( n19739 , n15252 , n6027 );
    nor g12548 ( n29052 , n12379 , n17488 );
    or g12549 ( n2320 , n22634 , n25709 );
    or g12550 ( n3520 , n6964 , n29828 );
    not g12551 ( n1945 , n24014 );
    nor g12552 ( n20746 , n28075 , n7880 );
    xnor g12553 ( n31892 , n8237 , n5703 );
    or g12554 ( n22727 , n24118 , n11698 );
    and g12555 ( n22707 , n29483 , n21241 );
    not g12556 ( n18989 , n23182 );
    not g12557 ( n18816 , n14445 );
    or g12558 ( n8537 , n27434 , n20516 );
    xnor g12559 ( n21418 , n9830 , n11294 );
    not g12560 ( n29829 , n5709 );
    not g12561 ( n25212 , n27559 );
    xnor g12562 ( n13114 , n13178 , n22586 );
    or g12563 ( n30361 , n3387 , n5105 );
    buf g12564 ( n24266 , n19976 );
    not g12565 ( n31956 , n13084 );
    xnor g12566 ( n8370 , n28397 , n2925 );
    and g12567 ( n26074 , n400 , n20869 );
    or g12568 ( n9175 , n12664 , n11028 );
    not g12569 ( n13419 , n7701 );
    xnor g12570 ( n1382 , n1592 , n12481 );
    not g12571 ( n23259 , n1813 );
    xnor g12572 ( n9391 , n3183 , n15141 );
    not g12573 ( n18333 , n20434 );
    not g12574 ( n29332 , n30303 );
    xnor g12575 ( n28261 , n26961 , n10433 );
    not g12576 ( n18587 , n30438 );
    or g12577 ( n23005 , n22678 , n29060 );
    or g12578 ( n5084 , n5955 , n24220 );
    xnor g12579 ( n23199 , n2002 , n22281 );
    and g12580 ( n16557 , n9242 , n8009 );
    nor g12581 ( n18249 , n28825 , n6253 );
    or g12582 ( n12650 , n20236 , n25997 );
    and g12583 ( n16915 , n26965 , n17787 );
    not g12584 ( n856 , n2529 );
    xnor g12585 ( n25515 , n31838 , n23936 );
    or g12586 ( n7178 , n25203 , n28707 );
    xnor g12587 ( n15619 , n9648 , n6204 );
    or g12588 ( n211 , n15799 , n5152 );
    or g12589 ( n14722 , n6062 , n27944 );
    not g12590 ( n11600 , n5511 );
    not g12591 ( n23209 , n30158 );
    xnor g12592 ( n25568 , n340 , n21986 );
    xnor g12593 ( n11267 , n31401 , n3641 );
    xnor g12594 ( n11775 , n137 , n27704 );
    and g12595 ( n17683 , n12925 , n8552 );
    and g12596 ( n5509 , n15903 , n24419 );
    and g12597 ( n8489 , n3268 , n25760 );
    xnor g12598 ( n2398 , n1299 , n13888 );
    nor g12599 ( n2108 , n8577 , n29252 );
    and g12600 ( n2239 , n11882 , n23036 );
    xnor g12601 ( n19970 , n15710 , n26151 );
    nor g12602 ( n8753 , n27787 , n11415 );
    xnor g12603 ( n5088 , n26835 , n16010 );
    not g12604 ( n25492 , n28845 );
    or g12605 ( n10744 , n30908 , n13680 );
    xnor g12606 ( n16271 , n30715 , n13962 );
    nor g12607 ( n13206 , n15652 , n19353 );
    or g12608 ( n19416 , n13517 , n20456 );
    not g12609 ( n13006 , n3101 );
    xnor g12610 ( n11636 , n25287 , n22848 );
    and g12611 ( n8695 , n22183 , n21517 );
    not g12612 ( n1950 , n12680 );
    not g12613 ( n372 , n13659 );
    xor g12614 ( n20708 , n27834 , n22677 );
    not g12615 ( n21039 , n26004 );
    nor g12616 ( n8731 , n13913 , n5110 );
    not g12617 ( n29162 , n30366 );
    xor g12618 ( n23976 , n17710 , n18551 );
    not g12619 ( n12344 , n4851 );
    or g12620 ( n13327 , n30275 , n12221 );
    not g12621 ( n5800 , n18869 );
    or g12622 ( n15136 , n22151 , n2324 );
    and g12623 ( n5932 , n6299 , n29997 );
    not g12624 ( n11450 , n30331 );
    and g12625 ( n12350 , n13202 , n12334 );
    not g12626 ( n15965 , n5498 );
    and g12627 ( n29533 , n10173 , n18405 );
    not g12628 ( n18078 , n6655 );
    and g12629 ( n21416 , n9761 , n6185 );
    nor g12630 ( n23728 , n31120 , n25364 );
    and g12631 ( n4091 , n6825 , n28189 );
    not g12632 ( n3536 , n9301 );
    not g12633 ( n27348 , n31100 );
    xnor g12634 ( n14166 , n9041 , n18959 );
    xnor g12635 ( n19222 , n18207 , n16406 );
    xnor g12636 ( n23401 , n20855 , n20224 );
    xor g12637 ( n7064 , n939 , n2757 );
    or g12638 ( n9767 , n4669 , n25812 );
    not g12639 ( n26941 , n30690 );
    not g12640 ( n28471 , n807 );
    not g12641 ( n28027 , n8761 );
    xnor g12642 ( n7904 , n13483 , n22341 );
    xnor g12643 ( n20900 , n11626 , n4990 );
    xnor g12644 ( n13059 , n25604 , n27660 );
    xnor g12645 ( n15744 , n9187 , n17995 );
    or g12646 ( n11642 , n18612 , n5111 );
    or g12647 ( n24791 , n6715 , n25404 );
    buf g12648 ( n26581 , n20914 );
    or g12649 ( n22229 , n10727 , n30324 );
    xnor g12650 ( n10031 , n30245 , n23770 );
    or g12651 ( n1851 , n21270 , n13606 );
    or g12652 ( n29241 , n23726 , n31119 );
    nor g12653 ( n28731 , n27632 , n27330 );
    and g12654 ( n2786 , n743 , n27890 );
    xnor g12655 ( n16233 , n12644 , n29194 );
    xnor g12656 ( n5390 , n10735 , n20641 );
    nor g12657 ( n17789 , n8701 , n16536 );
    xnor g12658 ( n4773 , n15200 , n2006 );
    and g12659 ( n11774 , n21991 , n5177 );
    not g12660 ( n8758 , n19467 );
    or g12661 ( n19391 , n28087 , n10931 );
    not g12662 ( n12652 , n12073 );
    xnor g12663 ( n30294 , n6264 , n16932 );
    xnor g12664 ( n10689 , n14327 , n16825 );
    not g12665 ( n4907 , n15145 );
    or g12666 ( n23939 , n26992 , n4110 );
    not g12667 ( n9711 , n7980 );
    nor g12668 ( n1015 , n15161 , n1306 );
    and g12669 ( n22761 , n25713 , n31666 );
    not g12670 ( n7625 , n14961 );
    or g12671 ( n17420 , n26205 , n6990 );
    or g12672 ( n22663 , n19941 , n25226 );
    and g12673 ( n5687 , n30813 , n12959 );
    xnor g12674 ( n9427 , n6484 , n738 );
    xnor g12675 ( n21071 , n11525 , n18729 );
    xnor g12676 ( n5998 , n2378 , n16299 );
    not g12677 ( n10261 , n13006 );
    not g12678 ( n23241 , n22618 );
    xnor g12679 ( n18943 , n6000 , n548 );
    or g12680 ( n7702 , n29606 , n7117 );
    not g12681 ( n10558 , n24940 );
    not g12682 ( n29975 , n27883 );
    and g12683 ( n2641 , n24211 , n30509 );
    and g12684 ( n19275 , n2002 , n26216 );
    not g12685 ( n10969 , n27075 );
    not g12686 ( n15410 , n5839 );
    xnor g12687 ( n7743 , n12355 , n17090 );
    and g12688 ( n26281 , n30668 , n28177 );
    xnor g12689 ( n12838 , n11454 , n2167 );
    or g12690 ( n27451 , n13643 , n32032 );
    not g12691 ( n24275 , n14195 );
    not g12692 ( n12075 , n17756 );
    not g12693 ( n6551 , n9414 );
    or g12694 ( n3777 , n29184 , n967 );
    not g12695 ( n3702 , n31519 );
    or g12696 ( n18270 , n956 , n3642 );
    xnor g12697 ( n23938 , n18253 , n22075 );
    not g12698 ( n29759 , n3726 );
    not g12699 ( n19366 , n9358 );
    and g12700 ( n3872 , n5372 , n21776 );
    or g12701 ( n14678 , n10647 , n18857 );
    or g12702 ( n27464 , n12636 , n21164 );
    xnor g12703 ( n132 , n16235 , n20039 );
    xnor g12704 ( n28160 , n17959 , n12871 );
    or g12705 ( n28556 , n22316 , n21606 );
    not g12706 ( n1344 , n29733 );
    nor g12707 ( n149 , n19720 , n26825 );
    xnor g12708 ( n29941 , n25941 , n21250 );
    nor g12709 ( n23718 , n15516 , n31443 );
    not g12710 ( n3898 , n24608 );
    xnor g12711 ( n9367 , n29081 , n2163 );
    not g12712 ( n28791 , n22232 );
    or g12713 ( n13696 , n14659 , n8465 );
    xnor g12714 ( n24260 , n2925 , n1095 );
    or g12715 ( n28361 , n846 , n19690 );
    or g12716 ( n27999 , n11479 , n18461 );
    not g12717 ( n3140 , n228 );
    nor g12718 ( n14078 , n30411 , n26082 );
    or g12719 ( n3328 , n20442 , n27724 );
    not g12720 ( n28617 , n3405 );
    not g12721 ( n12140 , n7354 );
    xnor g12722 ( n13275 , n26140 , n554 );
    xnor g12723 ( n11178 , n4463 , n24874 );
    and g12724 ( n19842 , n19646 , n27043 );
    or g12725 ( n6288 , n9571 , n19166 );
    nor g12726 ( n8331 , n17496 , n24961 );
    or g12727 ( n20478 , n6130 , n30200 );
    xnor g12728 ( n6 , n7629 , n27048 );
    nor g12729 ( n25014 , n21896 , n2537 );
    not g12730 ( n3005 , n5299 );
    or g12731 ( n19301 , n7728 , n18853 );
    not g12732 ( n7690 , n25858 );
    xnor g12733 ( n19241 , n24239 , n22958 );
    not g12734 ( n11671 , n30801 );
    and g12735 ( n3178 , n30708 , n5639 );
    and g12736 ( n16167 , n14762 , n13456 );
    and g12737 ( n13316 , n15621 , n6203 );
    or g12738 ( n18476 , n30779 , n28924 );
    or g12739 ( n8102 , n27488 , n20935 );
    xor g12740 ( n31682 , n18586 , n2866 );
    and g12741 ( n5326 , n15304 , n18638 );
    not g12742 ( n27205 , n27162 );
    not g12743 ( n22442 , n29807 );
    not g12744 ( n4435 , n21198 );
    or g12745 ( n22805 , n9015 , n3667 );
    not g12746 ( n14715 , n2264 );
    and g12747 ( n18659 , n14866 , n24960 );
    and g12748 ( n3159 , n9755 , n25356 );
    xnor g12749 ( n6905 , n15653 , n22237 );
    not g12750 ( n10202 , n2217 );
    or g12751 ( n8432 , n3037 , n10969 );
    not g12752 ( n17236 , n2700 );
    xnor g12753 ( n26859 , n6134 , n26479 );
    or g12754 ( n20614 , n6360 , n29592 );
    and g12755 ( n27241 , n27967 , n19720 );
    not g12756 ( n13879 , n10146 );
    not g12757 ( n25063 , n23960 );
    or g12758 ( n31488 , n30765 , n22725 );
    xnor g12759 ( n14401 , n22393 , n107 );
    xnor g12760 ( n16438 , n20492 , n7017 );
    xnor g12761 ( n10024 , n5691 , n7622 );
    xnor g12762 ( n7234 , n8127 , n8922 );
    and g12763 ( n6523 , n30208 , n27832 );
    or g12764 ( n8588 , n1895 , n9199 );
    or g12765 ( n18079 , n16733 , n13347 );
    xnor g12766 ( n23741 , n22490 , n31855 );
    or g12767 ( n14664 , n29705 , n9391 );
    and g12768 ( n31041 , n21959 , n3165 );
    xnor g12769 ( n2179 , n12998 , n24988 );
    and g12770 ( n24492 , n27306 , n16293 );
    xnor g12771 ( n6636 , n5162 , n27033 );
    xnor g12772 ( n18300 , n29002 , n11541 );
    xnor g12773 ( n15220 , n15836 , n24369 );
    not g12774 ( n23327 , n780 );
    xnor g12775 ( n365 , n22959 , n28115 );
    not g12776 ( n23811 , n23998 );
    nor g12777 ( n9267 , n13725 , n16357 );
    or g12778 ( n11129 , n26395 , n5599 );
    not g12779 ( n1551 , n10114 );
    nor g12780 ( n19764 , n3936 , n30904 );
    and g12781 ( n14461 , n2402 , n98 );
    xnor g12782 ( n5103 , n25413 , n7676 );
    not g12783 ( n7335 , n17305 );
    or g12784 ( n15811 , n2898 , n7381 );
    not g12785 ( n23510 , n8057 );
    nor g12786 ( n13050 , n29296 , n28630 );
    xnor g12787 ( n31012 , n23315 , n19670 );
    not g12788 ( n20987 , n19187 );
    not g12789 ( n15290 , n20435 );
    xnor g12790 ( n23430 , n7681 , n8762 );
    xnor g12791 ( n4439 , n10715 , n7492 );
    not g12792 ( n6181 , n14477 );
    or g12793 ( n8276 , n10856 , n3872 );
    and g12794 ( n15478 , n21623 , n9867 );
    nor g12795 ( n11067 , n27501 , n26661 );
    and g12796 ( n6881 , n29506 , n28127 );
    xnor g12797 ( n30648 , n21485 , n23232 );
    xnor g12798 ( n15024 , n28544 , n6647 );
    not g12799 ( n5435 , n6365 );
    xnor g12800 ( n19855 , n18143 , n5873 );
    or g12801 ( n23450 , n350 , n18990 );
    xnor g12802 ( n21322 , n6665 , n20885 );
    or g12803 ( n27688 , n1518 , n25275 );
    xnor g12804 ( n17918 , n436 , n22500 );
    and g12805 ( n7228 , n31318 , n823 );
    xnor g12806 ( n6687 , n6589 , n2129 );
    and g12807 ( n22286 , n14405 , n1535 );
    or g12808 ( n6714 , n14690 , n29440 );
    or g12809 ( n2692 , n5861 , n15246 );
    and g12810 ( n26157 , n9012 , n29463 );
    or g12811 ( n271 , n23312 , n21116 );
    nor g12812 ( n16475 , n30744 , n29929 );
    xnor g12813 ( n21716 , n438 , n4280 );
    nor g12814 ( n6584 , n27922 , n7242 );
    not g12815 ( n30927 , n12325 );
    or g12816 ( n31541 , n16605 , n10399 );
    nor g12817 ( n15989 , n9039 , n18283 );
    or g12818 ( n670 , n27684 , n25187 );
    not g12819 ( n26083 , n20704 );
    and g12820 ( n14494 , n5347 , n30738 );
    or g12821 ( n2580 , n12657 , n24729 );
    xor g12822 ( n16932 , n10862 , n13859 );
    not g12823 ( n15930 , n29708 );
    nor g12824 ( n12744 , n15842 , n2358 );
    or g12825 ( n25894 , n26867 , n14828 );
    not g12826 ( n20544 , n17575 );
    not g12827 ( n17424 , n18161 );
    not g12828 ( n9682 , n22778 );
    not g12829 ( n23834 , n18060 );
    xnor g12830 ( n11252 , n28638 , n3782 );
    not g12831 ( n28741 , n28431 );
    and g12832 ( n2 , n8951 , n28582 );
    xnor g12833 ( n17104 , n7410 , n16686 );
    not g12834 ( n4629 , n14967 );
    not g12835 ( n15309 , n9681 );
    not g12836 ( n27770 , n22280 );
    not g12837 ( n8667 , n31160 );
    and g12838 ( n8287 , n30747 , n29548 );
    xnor g12839 ( n24217 , n22343 , n10914 );
    xnor g12840 ( n4171 , n9098 , n18307 );
    not g12841 ( n666 , n31575 );
    not g12842 ( n30817 , n28252 );
    xnor g12843 ( n11343 , n4339 , n3641 );
    and g12844 ( n2565 , n6386 , n19695 );
    nor g12845 ( n24903 , n1113 , n8791 );
    or g12846 ( n26172 , n25698 , n2364 );
    xnor g12847 ( n24258 , n24169 , n23937 );
    or g12848 ( n3054 , n27133 , n10574 );
    nor g12849 ( n27286 , n20799 , n25902 );
    or g12850 ( n5508 , n1720 , n12001 );
    nor g12851 ( n28525 , n8736 , n9716 );
    or g12852 ( n20547 , n24552 , n25174 );
    xnor g12853 ( n536 , n25656 , n296 );
    nor g12854 ( n15583 , n30268 , n7687 );
    or g12855 ( n8633 , n5892 , n14236 );
    not g12856 ( n3039 , n29249 );
    xnor g12857 ( n22022 , n26000 , n10456 );
    not g12858 ( n1640 , n4393 );
    not g12859 ( n12429 , n25284 );
    or g12860 ( n114 , n29293 , n9337 );
    xnor g12861 ( n1445 , n23316 , n8385 );
    and g12862 ( n18099 , n25822 , n25998 );
    not g12863 ( n7199 , n29002 );
    not g12864 ( n30790 , n24990 );
    not g12865 ( n16304 , n358 );
    not g12866 ( n29756 , n2781 );
    and g12867 ( n8932 , n2896 , n15359 );
    not g12868 ( n9718 , n27364 );
    not g12869 ( n31074 , n19405 );
    or g12870 ( n2930 , n20967 , n4117 );
    or g12871 ( n24971 , n12666 , n29027 );
    xnor g12872 ( n28707 , n14101 , n24206 );
    xnor g12873 ( n21659 , n25405 , n22349 );
    and g12874 ( n12810 , n29134 , n27591 );
    and g12875 ( n24954 , n20911 , n31071 );
    nor g12876 ( n29291 , n664 , n29249 );
    not g12877 ( n10237 , n21122 );
    and g12878 ( n15031 , n6854 , n2293 );
    and g12879 ( n14778 , n8494 , n22283 );
    xnor g12880 ( n26676 , n25542 , n29832 );
    or g12881 ( n14953 , n16528 , n7494 );
    or g12882 ( n6561 , n24540 , n19752 );
    and g12883 ( n21048 , n18261 , n19129 );
    not g12884 ( n4678 , n31193 );
    and g12885 ( n1211 , n27138 , n13324 );
    or g12886 ( n17049 , n19936 , n17372 );
    or g12887 ( n14179 , n27054 , n29924 );
    not g12888 ( n5265 , n10083 );
    xnor g12889 ( n2828 , n3637 , n27058 );
    not g12890 ( n15892 , n24620 );
    and g12891 ( n8888 , n27718 , n4050 );
    and g12892 ( n26952 , n27337 , n12247 );
    xnor g12893 ( n25470 , n23130 , n14769 );
    or g12894 ( n13202 , n25861 , n23690 );
    not g12895 ( n1831 , n8758 );
    and g12896 ( n15415 , n22839 , n10953 );
    not g12897 ( n4491 , n25318 );
    not g12898 ( n847 , n19928 );
    not g12899 ( n788 , n18599 );
    not g12900 ( n3484 , n6036 );
    not g12901 ( n24166 , n22166 );
    nor g12902 ( n5425 , n17588 , n9407 );
    or g12903 ( n26050 , n22612 , n28751 );
    not g12904 ( n8910 , n13283 );
    not g12905 ( n3604 , n8964 );
    xnor g12906 ( n29623 , n23785 , n5085 );
    or g12907 ( n26135 , n3307 , n30744 );
    or g12908 ( n4389 , n6233 , n11936 );
    or g12909 ( n25321 , n16185 , n20893 );
    or g12910 ( n7828 , n14721 , n28481 );
    not g12911 ( n6456 , n31066 );
    xor g12912 ( n22295 , n114 , n31094 );
    nor g12913 ( n26098 , n20620 , n24854 );
    xnor g12914 ( n5446 , n3885 , n28940 );
    or g12915 ( n13173 , n16284 , n17597 );
    xnor g12916 ( n16578 , n11784 , n21349 );
    and g12917 ( n11673 , n19900 , n29887 );
    xnor g12918 ( n13309 , n22951 , n5258 );
    xnor g12919 ( n21161 , n30283 , n27565 );
    not g12920 ( n6347 , n24356 );
    xnor g12921 ( n15060 , n12919 , n32027 );
    or g12922 ( n23191 , n7714 , n18860 );
    xnor g12923 ( n26285 , n16098 , n29759 );
    xnor g12924 ( n26799 , n29696 , n3921 );
    or g12925 ( n16876 , n22401 , n14932 );
    not g12926 ( n17063 , n11526 );
    or g12927 ( n20376 , n17807 , n8044 );
    not g12928 ( n22646 , n31168 );
    not g12929 ( n18921 , n14994 );
    and g12930 ( n369 , n21730 , n22737 );
    xnor g12931 ( n22799 , n3477 , n17249 );
    nor g12932 ( n22558 , n20525 , n11178 );
    nor g12933 ( n16509 , n22886 , n28689 );
    or g12934 ( n457 , n8917 , n12989 );
    not g12935 ( n25814 , n5765 );
    not g12936 ( n1479 , n10793 );
    xnor g12937 ( n28773 , n4890 , n11127 );
    and g12938 ( n23760 , n20123 , n855 );
    nor g12939 ( n8306 , n7214 , n18119 );
    and g12940 ( n5436 , n6453 , n12373 );
    xnor g12941 ( n15283 , n13128 , n21889 );
    xnor g12942 ( n31166 , n4069 , n19317 );
    not g12943 ( n311 , n26833 );
    not g12944 ( n21167 , n6661 );
    not g12945 ( n26601 , n12409 );
    and g12946 ( n10740 , n13532 , n23480 );
    not g12947 ( n18242 , n8210 );
    not g12948 ( n20293 , n16209 );
    not g12949 ( n22712 , n14368 );
    or g12950 ( n31870 , n20762 , n20405 );
    or g12951 ( n4797 , n30201 , n1422 );
    not g12952 ( n19953 , n11132 );
    and g12953 ( n20915 , n5824 , n25683 );
    or g12954 ( n8691 , n10803 , n83 );
    nor g12955 ( n1306 , n11230 , n28396 );
    not g12956 ( n29163 , n15362 );
    not g12957 ( n20350 , n828 );
    and g12958 ( n22483 , n4230 , n22898 );
    not g12959 ( n23648 , n11838 );
    and g12960 ( n10592 , n8795 , n8254 );
    xnor g12961 ( n24549 , n10116 , n16993 );
    nor g12962 ( n6508 , n31228 , n27512 );
    nor g12963 ( n24830 , n24302 , n31956 );
    or g12964 ( n12606 , n28039 , n13248 );
    not g12965 ( n11497 , n21963 );
    nor g12966 ( n17116 , n18198 , n9445 );
    not g12967 ( n6267 , n30122 );
    xnor g12968 ( n17234 , n11394 , n802 );
    or g12969 ( n14068 , n2178 , n6092 );
    xnor g12970 ( n27621 , n26733 , n24622 );
    and g12971 ( n14637 , n29579 , n791 );
    xnor g12972 ( n15940 , n4798 , n4169 );
    and g12973 ( n3348 , n28455 , n15688 );
    not g12974 ( n5539 , n4567 );
    or g12975 ( n20622 , n13271 , n14228 );
    and g12976 ( n24000 , n9127 , n11087 );
    or g12977 ( n16814 , n28517 , n12469 );
    not g12978 ( n23541 , n6650 );
    or g12979 ( n14059 , n7860 , n20990 );
    or g12980 ( n45 , n2854 , n13483 );
    and g12981 ( n7806 , n26421 , n23753 );
    or g12982 ( n26126 , n22578 , n6269 );
    or g12983 ( n28123 , n17601 , n21730 );
    not g12984 ( n3519 , n20249 );
    or g12985 ( n23347 , n28355 , n6763 );
    not g12986 ( n2571 , n22549 );
    xnor g12987 ( n9361 , n14010 , n5462 );
    and g12988 ( n75 , n24078 , n11794 );
    not g12989 ( n5631 , n84 );
    and g12990 ( n15065 , n712 , n2265 );
    or g12991 ( n6536 , n11372 , n21714 );
    xnor g12992 ( n5148 , n14872 , n6249 );
    and g12993 ( n6263 , n10878 , n4553 );
    not g12994 ( n10962 , n30504 );
    or g12995 ( n18982 , n22635 , n20953 );
    not g12996 ( n20476 , n22717 );
    xnor g12997 ( n26248 , n27732 , n29415 );
    or g12998 ( n28461 , n6246 , n30238 );
    and g12999 ( n26578 , n11365 , n29123 );
    or g13000 ( n20314 , n5563 , n7307 );
    not g13001 ( n20742 , n15764 );
    buf g13002 ( n18496 , n19902 );
    or g13003 ( n1779 , n18338 , n12137 );
    xnor g13004 ( n21192 , n10927 , n18794 );
    or g13005 ( n8720 , n11360 , n2814 );
    and g13006 ( n22485 , n552 , n21874 );
    or g13007 ( n12296 , n20956 , n31024 );
    not g13008 ( n27668 , n12080 );
    and g13009 ( n17552 , n11825 , n26614 );
    not g13010 ( n7740 , n7161 );
    and g13011 ( n5279 , n24188 , n27202 );
    xnor g13012 ( n27368 , n30055 , n22801 );
    not g13013 ( n4198 , n4087 );
    and g13014 ( n8895 , n21155 , n31716 );
    not g13015 ( n5294 , n9485 );
    and g13016 ( n19773 , n6046 , n8418 );
    or g13017 ( n219 , n28260 , n25072 );
    xnor g13018 ( n24797 , n18662 , n28781 );
    not g13019 ( n27154 , n13356 );
    xnor g13020 ( n2649 , n24837 , n23115 );
    not g13021 ( n3498 , n30195 );
    xnor g13022 ( n16718 , n18261 , n3817 );
    nor g13023 ( n6529 , n20905 , n11416 );
    or g13024 ( n20513 , n22474 , n13458 );
    not g13025 ( n8284 , n18695 );
    or g13026 ( n25129 , n24202 , n15056 );
    not g13027 ( n27873 , n4335 );
    or g13028 ( n22495 , n7024 , n27899 );
    and g13029 ( n28481 , n18756 , n26417 );
    xnor g13030 ( n8427 , n19300 , n30514 );
    xnor g13031 ( n7107 , n14354 , n260 );
    xnor g13032 ( n26966 , n14296 , n18379 );
    and g13033 ( n13566 , n17716 , n6482 );
    or g13034 ( n9454 , n7776 , n21059 );
    xnor g13035 ( n12488 , n19812 , n15521 );
    not g13036 ( n24063 , n15045 );
    and g13037 ( n19724 , n8224 , n10568 );
    xnor g13038 ( n27243 , n13002 , n10709 );
    xnor g13039 ( n28957 , n11551 , n22460 );
    or g13040 ( n24278 , n5392 , n31289 );
    or g13041 ( n20886 , n14094 , n27617 );
    and g13042 ( n13670 , n3008 , n17267 );
    xnor g13043 ( n16402 , n3062 , n5374 );
    nor g13044 ( n18018 , n2985 , n16872 );
    xnor g13045 ( n30323 , n1799 , n115 );
    and g13046 ( n7467 , n16644 , n30280 );
    not g13047 ( n11803 , n4656 );
    and g13048 ( n8091 , n586 , n29765 );
    nor g13049 ( n14764 , n13616 , n13945 );
    not g13050 ( n4910 , n16420 );
    not g13051 ( n31707 , n26963 );
    not g13052 ( n7280 , n16111 );
    xnor g13053 ( n13500 , n16832 , n18589 );
    xor g13054 ( n31436 , n12631 , n2353 );
    not g13055 ( n25245 , n12564 );
    and g13056 ( n29110 , n25333 , n3321 );
    and g13057 ( n23257 , n2145 , n25653 );
    or g13058 ( n5875 , n18554 , n25348 );
    not g13059 ( n7224 , n10497 );
    or g13060 ( n25607 , n13820 , n16211 );
    or g13061 ( n21721 , n17655 , n25229 );
    not g13062 ( n19951 , n11861 );
    xnor g13063 ( n22159 , n30728 , n10451 );
    and g13064 ( n3881 , n12927 , n20241 );
    not g13065 ( n17974 , n21774 );
    xnor g13066 ( n27088 , n22942 , n5300 );
    or g13067 ( n22883 , n4477 , n5216 );
    xnor g13068 ( n25966 , n28368 , n29239 );
    not g13069 ( n19988 , n14288 );
    not g13070 ( n16313 , n14834 );
    or g13071 ( n245 , n4531 , n6240 );
    xnor g13072 ( n23167 , n17429 , n31481 );
    nor g13073 ( n10806 , n2684 , n1218 );
    not g13074 ( n15717 , n8338 );
    xor g13075 ( n12687 , n25435 , n4092 );
    or g13076 ( n26363 , n17523 , n9107 );
    or g13077 ( n20073 , n4449 , n23385 );
    and g13078 ( n17976 , n28317 , n31587 );
    or g13079 ( n16622 , n27470 , n31048 );
    or g13080 ( n9292 , n29036 , n21998 );
    xnor g13081 ( n8949 , n22729 , n745 );
    nor g13082 ( n29517 , n5348 , n14317 );
    or g13083 ( n13063 , n28433 , n14035 );
    not g13084 ( n18166 , n31078 );
    nor g13085 ( n15138 , n23518 , n302 );
    not g13086 ( n23736 , n20815 );
    and g13087 ( n30442 , n3320 , n9511 );
    or g13088 ( n6008 , n21086 , n696 );
    not g13089 ( n12952 , n21771 );
    xnor g13090 ( n17119 , n22043 , n10841 );
    xnor g13091 ( n3676 , n18790 , n26987 );
    xor g13092 ( n4090 , n8864 , n3844 );
    xnor g13093 ( n3510 , n4656 , n24118 );
    and g13094 ( n13946 , n28446 , n23457 );
    or g13095 ( n31820 , n24064 , n31931 );
    not g13096 ( n708 , n27435 );
    and g13097 ( n7493 , n30338 , n18781 );
    or g13098 ( n4063 , n19654 , n18980 );
    not g13099 ( n22082 , n16392 );
    xnor g13100 ( n30909 , n8397 , n12857 );
    or g13101 ( n20640 , n10691 , n5889 );
    or g13102 ( n13784 , n735 , n11012 );
    nor g13103 ( n13694 , n29138 , n21106 );
    and g13104 ( n21586 , n8746 , n10035 );
    xnor g13105 ( n20909 , n26793 , n9220 );
    xnor g13106 ( n12975 , n7442 , n4698 );
    xnor g13107 ( n27361 , n19906 , n7059 );
    not g13108 ( n24468 , n13265 );
    not g13109 ( n31072 , n1494 );
    and g13110 ( n31495 , n24529 , n19320 );
    xnor g13111 ( n14015 , n15048 , n9922 );
    xnor g13112 ( n11100 , n21501 , n26242 );
    and g13113 ( n4643 , n18742 , n23950 );
    not g13114 ( n31462 , n6394 );
    nor g13115 ( n18051 , n14040 , n25403 );
    and g13116 ( n22732 , n17434 , n6536 );
    not g13117 ( n30301 , n30593 );
    not g13118 ( n19218 , n7891 );
    xnor g13119 ( n18915 , n408 , n21272 );
    or g13120 ( n7049 , n1670 , n30923 );
    not g13121 ( n29071 , n11869 );
    and g13122 ( n21171 , n6671 , n30012 );
    or g13123 ( n12115 , n28874 , n17544 );
    and g13124 ( n22288 , n22000 , n21965 );
    xnor g13125 ( n12788 , n767 , n6939 );
    and g13126 ( n22481 , n25542 , n31235 );
    not g13127 ( n2694 , n21653 );
    xnor g13128 ( n19309 , n9310 , n4662 );
    not g13129 ( n27026 , n1720 );
    xnor g13130 ( n6950 , n25814 , n6163 );
    not g13131 ( n25278 , n31501 );
    not g13132 ( n21049 , n28807 );
    not g13133 ( n8186 , n20543 );
    xnor g13134 ( n8095 , n23751 , n22716 );
    xor g13135 ( n2422 , n12292 , n17281 );
    or g13136 ( n27494 , n20041 , n20793 );
    and g13137 ( n7368 , n23528 , n18170 );
    or g13138 ( n7406 , n12763 , n6921 );
    and g13139 ( n9110 , n14244 , n9493 );
    not g13140 ( n30863 , n31182 );
    or g13141 ( n14541 , n30135 , n30445 );
    or g13142 ( n25787 , n4306 , n15106 );
    not g13143 ( n23705 , n22423 );
    xnor g13144 ( n27537 , n24370 , n2451 );
    not g13145 ( n17356 , n18502 );
    xnor g13146 ( n12816 , n19506 , n11612 );
    not g13147 ( n1114 , n11982 );
    not g13148 ( n26560 , n5133 );
    xnor g13149 ( n4983 , n27437 , n12297 );
    not g13150 ( n4145 , n19839 );
    xnor g13151 ( n29538 , n12390 , n21259 );
    xnor g13152 ( n13528 , n13311 , n4925 );
    not g13153 ( n16230 , n22316 );
    and g13154 ( n21527 , n8196 , n21280 );
    not g13155 ( n933 , n3861 );
    not g13156 ( n17338 , n19597 );
    or g13157 ( n21319 , n19074 , n1338 );
    not g13158 ( n7111 , n2388 );
    not g13159 ( n21677 , n13158 );
    and g13160 ( n6571 , n30436 , n13719 );
    or g13161 ( n31938 , n7400 , n29728 );
    xnor g13162 ( n6931 , n30287 , n9336 );
    not g13163 ( n14946 , n2339 );
    xnor g13164 ( n24291 , n3764 , n9935 );
    or g13165 ( n605 , n18583 , n13602 );
    not g13166 ( n30396 , n11468 );
    xnor g13167 ( n16498 , n9576 , n14095 );
    not g13168 ( n28106 , n14241 );
    xnor g13169 ( n3665 , n14451 , n30529 );
    xnor g13170 ( n29418 , n25725 , n13920 );
    not g13171 ( n2461 , n2268 );
    not g13172 ( n17820 , n4361 );
    or g13173 ( n8564 , n9228 , n22451 );
    not g13174 ( n5075 , n7284 );
    not g13175 ( n20890 , n14657 );
    xnor g13176 ( n30722 , n13817 , n16132 );
    xnor g13177 ( n21521 , n23176 , n30196 );
    not g13178 ( n7396 , n19976 );
    not g13179 ( n19692 , n26636 );
    xor g13180 ( n11738 , n26626 , n15 );
    or g13181 ( n9329 , n15607 , n8034 );
    or g13182 ( n30598 , n6186 , n29068 );
    not g13183 ( n22581 , n12779 );
    or g13184 ( n30511 , n2624 , n21857 );
    xnor g13185 ( n25498 , n20233 , n27453 );
    xnor g13186 ( n6110 , n26512 , n3034 );
    not g13187 ( n2668 , n18731 );
    not g13188 ( n22496 , n6217 );
    xnor g13189 ( n19548 , n6084 , n16873 );
    xnor g13190 ( n22205 , n16428 , n12154 );
    xnor g13191 ( n811 , n10320 , n22075 );
    and g13192 ( n26128 , n21596 , n7579 );
    not g13193 ( n23982 , n12056 );
    not g13194 ( n1145 , n4059 );
    xnor g13195 ( n16862 , n17078 , n31105 );
    or g13196 ( n25899 , n2280 , n20454 );
    xnor g13197 ( n25660 , n25697 , n20860 );
    xnor g13198 ( n23373 , n11658 , n7314 );
    xnor g13199 ( n29189 , n10033 , n7508 );
    not g13200 ( n31817 , n10220 );
    xnor g13201 ( n20006 , n13761 , n28502 );
    or g13202 ( n15197 , n320 , n7456 );
    and g13203 ( n4520 , n23031 , n5049 );
    or g13204 ( n22978 , n31727 , n6970 );
    nor g13205 ( n6042 , n2939 , n9877 );
    or g13206 ( n17160 , n27710 , n16687 );
    and g13207 ( n7062 , n30637 , n4835 );
    not g13208 ( n16884 , n22393 );
    or g13209 ( n29123 , n22643 , n23098 );
    or g13210 ( n20354 , n22268 , n27946 );
    not g13211 ( n23415 , n23476 );
    not g13212 ( n19437 , n2718 );
    not g13213 ( n13634 , n17190 );
    not g13214 ( n31677 , n20 );
    xnor g13215 ( n13547 , n739 , n32 );
    not g13216 ( n9803 , n7033 );
    xnor g13217 ( n30931 , n26753 , n5025 );
    not g13218 ( n8134 , n5118 );
    or g13219 ( n3561 , n18110 , n26273 );
    not g13220 ( n23519 , n28600 );
    xnor g13221 ( n24535 , n17483 , n22368 );
    and g13222 ( n22872 , n1164 , n26120 );
    xnor g13223 ( n27949 , n1635 , n3432 );
    xnor g13224 ( n14966 , n10949 , n13833 );
    not g13225 ( n20935 , n7839 );
    not g13226 ( n10641 , n22332 );
    nor g13227 ( n13991 , n15525 , n9783 );
    and g13228 ( n14771 , n641 , n4182 );
    xnor g13229 ( n24021 , n15236 , n27237 );
    and g13230 ( n7731 , n22028 , n763 );
    xnor g13231 ( n20836 , n19307 , n17822 );
    nor g13232 ( n7960 , n30245 , n12566 );
    not g13233 ( n8256 , n26920 );
    and g13234 ( n17544 , n27683 , n16136 );
    not g13235 ( n7246 , n10463 );
    or g13236 ( n20792 , n4605 , n16232 );
    not g13237 ( n30806 , n16831 );
    or g13238 ( n21756 , n20142 , n25437 );
    xnor g13239 ( n24682 , n5451 , n30831 );
    not g13240 ( n1477 , n8853 );
    not g13241 ( n29069 , n11920 );
    or g13242 ( n14748 , n23730 , n12133 );
    or g13243 ( n25746 , n6248 , n7567 );
    not g13244 ( n29881 , n15111 );
    xnor g13245 ( n3715 , n9604 , n24522 );
    or g13246 ( n4411 , n23181 , n29942 );
    xnor g13247 ( n17321 , n18567 , n24260 );
    xnor g13248 ( n17147 , n12986 , n21808 );
    xnor g13249 ( n20819 , n11646 , n6692 );
    and g13250 ( n12682 , n9149 , n24379 );
    or g13251 ( n6268 , n30141 , n21227 );
    xnor g13252 ( n14635 , n16604 , n29513 );
    xnor g13253 ( n24811 , n14406 , n23089 );
    and g13254 ( n24585 , n17490 , n30985 );
    not g13255 ( n15506 , n17748 );
    not g13256 ( n23433 , n6594 );
    xnor g13257 ( n17024 , n4475 , n5390 );
    xnor g13258 ( n4590 , n4678 , n13514 );
    nor g13259 ( n19661 , n17075 , n21323 );
    and g13260 ( n7295 , n25254 , n28441 );
    xnor g13261 ( n3234 , n19093 , n6141 );
    nor g13262 ( n4153 , n1828 , n10104 );
    or g13263 ( n19127 , n27824 , n28276 );
    not g13264 ( n31090 , n31584 );
    not g13265 ( n26853 , n6036 );
    nor g13266 ( n9299 , n31246 , n17123 );
    and g13267 ( n31402 , n28967 , n1625 );
    xnor g13268 ( n30056 , n30842 , n26401 );
    or g13269 ( n8756 , n2919 , n22539 );
    xnor g13270 ( n25467 , n4443 , n501 );
    not g13271 ( n787 , n25682 );
    and g13272 ( n27824 , n7344 , n19897 );
    nor g13273 ( n636 , n4179 , n26845 );
    or g13274 ( n7484 , n5189 , n14895 );
    xnor g13275 ( n5099 , n29679 , n22407 );
    and g13276 ( n11299 , n22193 , n3820 );
    or g13277 ( n28495 , n16069 , n174 );
    or g13278 ( n30782 , n717 , n5007 );
    nor g13279 ( n23896 , n20453 , n20823 );
    not g13280 ( n456 , n22691 );
    or g13281 ( n30613 , n14554 , n3539 );
    xnor g13282 ( n21405 , n27809 , n23697 );
    or g13283 ( n544 , n9591 , n73 );
    and g13284 ( n2487 , n29909 , n12367 );
    or g13285 ( n29379 , n22646 , n17090 );
    xnor g13286 ( n14091 , n22990 , n12356 );
    not g13287 ( n30586 , n22136 );
    xnor g13288 ( n31624 , n18611 , n20579 );
    not g13289 ( n17740 , n10364 );
    xnor g13290 ( n19505 , n27190 , n17591 );
    or g13291 ( n27545 , n9541 , n26651 );
    xnor g13292 ( n12352 , n15154 , n26888 );
    nor g13293 ( n11686 , n27962 , n23946 );
    not g13294 ( n8445 , n2106 );
    or g13295 ( n8606 , n16734 , n23718 );
    xnor g13296 ( n11187 , n6421 , n4702 );
    not g13297 ( n10092 , n17686 );
    not g13298 ( n2749 , n24857 );
    nor g13299 ( n24326 , n4310 , n30645 );
    xnor g13300 ( n2356 , n6155 , n15840 );
    not g13301 ( n22057 , n31526 );
    xnor g13302 ( n20594 , n12885 , n6512 );
    xnor g13303 ( n30114 , n1152 , n7760 );
    not g13304 ( n25994 , n28678 );
    or g13305 ( n28291 , n6398 , n9038 );
    nor g13306 ( n6601 , n5873 , n17561 );
    not g13307 ( n30398 , n9525 );
    xnor g13308 ( n18214 , n6197 , n5381 );
    not g13309 ( n7981 , n8890 );
    not g13310 ( n4615 , n23533 );
    xnor g13311 ( n122 , n3913 , n11257 );
    xnor g13312 ( n30954 , n1594 , n13480 );
    and g13313 ( n14572 , n7753 , n6842 );
    and g13314 ( n239 , n20875 , n27622 );
    or g13315 ( n14522 , n5870 , n13505 );
    not g13316 ( n5677 , n12998 );
    not g13317 ( n21044 , n29643 );
    xnor g13318 ( n10404 , n28554 , n28779 );
    not g13319 ( n30305 , n20607 );
    or g13320 ( n9148 , n28646 , n9961 );
    or g13321 ( n20230 , n29437 , n8971 );
    nor g13322 ( n11266 , n9080 , n6338 );
    not g13323 ( n29282 , n6565 );
    not g13324 ( n31745 , n6010 );
    xnor g13325 ( n23857 , n1183 , n4108 );
    nor g13326 ( n243 , n16449 , n6929 );
    xnor g13327 ( n26746 , n27933 , n17269 );
    and g13328 ( n25266 , n29275 , n23213 );
    and g13329 ( n14799 , n3852 , n12027 );
    xnor g13330 ( n26602 , n15215 , n2538 );
    nor g13331 ( n31770 , n7390 , n19196 );
    not g13332 ( n23266 , n27979 );
    not g13333 ( n24031 , n5718 );
    nor g13334 ( n27040 , n20667 , n28867 );
    not g13335 ( n2724 , n25510 );
    not g13336 ( n26731 , n974 );
    nor g13337 ( n28503 , n25708 , n25570 );
    or g13338 ( n11783 , n29826 , n13079 );
    not g13339 ( n20872 , n19704 );
    xnor g13340 ( n7389 , n8495 , n16090 );
    xnor g13341 ( n13049 , n4864 , n28058 );
    and g13342 ( n6761 , n29760 , n16346 );
    not g13343 ( n28066 , n16860 );
    nor g13344 ( n20122 , n27805 , n25982 );
    not g13345 ( n2574 , n26298 );
    and g13346 ( n29823 , n29233 , n3816 );
    xnor g13347 ( n11031 , n28816 , n15520 );
    or g13348 ( n13435 , n15500 , n25499 );
    or g13349 ( n15104 , n27299 , n8954 );
    not g13350 ( n14270 , n25690 );
    xnor g13351 ( n7033 , n22458 , n21552 );
    xnor g13352 ( n26462 , n13393 , n20632 );
    not g13353 ( n27 , n31191 );
    or g13354 ( n28775 , n19088 , n16042 );
    xnor g13355 ( n59 , n7305 , n21658 );
    xnor g13356 ( n13438 , n13391 , n7152 );
    xnor g13357 ( n24849 , n14661 , n10362 );
    and g13358 ( n10726 , n12085 , n3842 );
    nor g13359 ( n17846 , n8738 , n21840 );
    and g13360 ( n9018 , n3687 , n20741 );
    and g13361 ( n16025 , n18835 , n31311 );
    not g13362 ( n25535 , n20503 );
    xnor g13363 ( n17146 , n20231 , n24213 );
    or g13364 ( n19504 , n30771 , n24362 );
    xnor g13365 ( n8953 , n13136 , n4595 );
    not g13366 ( n23230 , n1867 );
    xnor g13367 ( n26593 , n4970 , n9057 );
    xnor g13368 ( n23838 , n6485 , n27469 );
    nor g13369 ( n30291 , n20069 , n5101 );
    xnor g13370 ( n16164 , n22444 , n16807 );
    xnor g13371 ( n2128 , n1193 , n13642 );
    and g13372 ( n21424 , n19938 , n14324 );
    xnor g13373 ( n19881 , n3259 , n6306 );
    and g13374 ( n12480 , n21319 , n15163 );
    nor g13375 ( n22192 , n10435 , n8392 );
    xnor g13376 ( n26830 , n21904 , n2109 );
    xnor g13377 ( n30910 , n18827 , n30029 );
    not g13378 ( n4994 , n29569 );
    or g13379 ( n29549 , n9235 , n11851 );
    not g13380 ( n16942 , n22867 );
    or g13381 ( n4635 , n10267 , n22462 );
    not g13382 ( n27132 , n13735 );
    xnor g13383 ( n27767 , n7763 , n13829 );
    and g13384 ( n14734 , n16627 , n31529 );
    not g13385 ( n18404 , n23079 );
    and g13386 ( n14174 , n13149 , n16238 );
    nor g13387 ( n29495 , n18002 , n30699 );
    and g13388 ( n24177 , n15798 , n23890 );
    or g13389 ( n262 , n31696 , n10271 );
    not g13390 ( n5240 , n23297 );
    nor g13391 ( n2371 , n5773 , n13664 );
    and g13392 ( n15602 , n6120 , n16546 );
    xnor g13393 ( n27427 , n11332 , n28192 );
    and g13394 ( n23610 , n21092 , n20287 );
    or g13395 ( n18213 , n9197 , n27821 );
    or g13396 ( n30762 , n21030 , n25135 );
    or g13397 ( n28153 , n13765 , n21050 );
    nor g13398 ( n19027 , n2308 , n19404 );
    or g13399 ( n2014 , n24670 , n29680 );
    or g13400 ( n24882 , n23883 , n29681 );
    xnor g13401 ( n18878 , n17200 , n22075 );
    or g13402 ( n28308 , n20285 , n8595 );
    nor g13403 ( n962 , n26396 , n17762 );
    not g13404 ( n18954 , n12200 );
    or g13405 ( n30619 , n8006 , n26452 );
    xnor g13406 ( n30707 , n9462 , n28474 );
    xnor g13407 ( n15077 , n21080 , n12857 );
    or g13408 ( n21511 , n12514 , n17455 );
    or g13409 ( n28522 , n16945 , n31533 );
    and g13410 ( n15864 , n2175 , n27161 );
    not g13411 ( n30479 , n7438 );
    nor g13412 ( n8261 , n9116 , n30601 );
    not g13413 ( n29774 , n29170 );
    and g13414 ( n15616 , n10824 , n13921 );
    xnor g13415 ( n27888 , n22129 , n23577 );
    or g13416 ( n10026 , n25886 , n6293 );
    not g13417 ( n1067 , n13602 );
    xnor g13418 ( n769 , n22845 , n18507 );
    not g13419 ( n13663 , n17141 );
    or g13420 ( n10371 , n27068 , n28902 );
    or g13421 ( n24742 , n5440 , n10473 );
    xnor g13422 ( n31696 , n28101 , n23987 );
    or g13423 ( n27817 , n5551 , n12166 );
    and g13424 ( n23393 , n28865 , n3923 );
    xnor g13425 ( n20782 , n29791 , n30351 );
    or g13426 ( n2637 , n445 , n16208 );
    xnor g13427 ( n20697 , n2925 , n3614 );
    or g13428 ( n14240 , n20957 , n5015 );
    nor g13429 ( n19945 , n4196 , n3269 );
    not g13430 ( n17915 , n27013 );
    xnor g13431 ( n6497 , n23585 , n21468 );
    and g13432 ( n6672 , n15160 , n8144 );
    and g13433 ( n20361 , n15817 , n4380 );
    and g13434 ( n19669 , n10023 , n7366 );
    and g13435 ( n13630 , n3790 , n23193 );
    xnor g13436 ( n7407 , n7354 , n8867 );
    not g13437 ( n18650 , n30697 );
    not g13438 ( n6199 , n2270 );
    and g13439 ( n2193 , n19253 , n27739 );
    xnor g13440 ( n5558 , n3353 , n8162 );
    or g13441 ( n30726 , n22350 , n28302 );
    or g13442 ( n18794 , n26910 , n24150 );
    xnor g13443 ( n18387 , n1935 , n16238 );
    not g13444 ( n5474 , n10947 );
    nor g13445 ( n21093 , n29414 , n6960 );
    or g13446 ( n21243 , n7014 , n28679 );
    and g13447 ( n18069 , n3851 , n31237 );
    or g13448 ( n20737 , n16516 , n22344 );
    xnor g13449 ( n7640 , n8311 , n2753 );
    or g13450 ( n7719 , n6948 , n18218 );
    or g13451 ( n14857 , n6540 , n15206 );
    or g13452 ( n3120 , n14174 , n13595 );
    not g13453 ( n11629 , n6475 );
    or g13454 ( n29853 , n2231 , n30733 );
    not g13455 ( n24547 , n5972 );
    or g13456 ( n9415 , n13412 , n18736 );
    not g13457 ( n10982 , n29437 );
    not g13458 ( n10639 , n18344 );
    not g13459 ( n1291 , n18155 );
    or g13460 ( n27096 , n23720 , n1033 );
    not g13461 ( n5438 , n24739 );
    xnor g13462 ( n24005 , n17820 , n26700 );
    xnor g13463 ( n22546 , n19784 , n22357 );
    not g13464 ( n23481 , n29756 );
    and g13465 ( n21378 , n19750 , n8684 );
    not g13466 ( n15677 , n7004 );
    nor g13467 ( n21150 , n13145 , n10982 );
    or g13468 ( n503 , n28511 , n27180 );
    not g13469 ( n28869 , n4847 );
    xnor g13470 ( n8422 , n22781 , n16417 );
    and g13471 ( n31335 , n28506 , n30973 );
    nor g13472 ( n21725 , n2231 , n3039 );
    or g13473 ( n11821 , n10750 , n11726 );
    or g13474 ( n29636 , n16005 , n19854 );
    not g13475 ( n3683 , n31128 );
    or g13476 ( n16506 , n12810 , n20502 );
    not g13477 ( n22005 , n23770 );
    or g13478 ( n22225 , n28156 , n7432 );
    and g13479 ( n10708 , n6878 , n4263 );
    not g13480 ( n26687 , n21277 );
    or g13481 ( n19070 , n11631 , n857 );
    and g13482 ( n28467 , n288 , n26641 );
    and g13483 ( n9787 , n13596 , n5720 );
    and g13484 ( n6333 , n14710 , n597 );
    xnor g13485 ( n15642 , n14640 , n28319 );
    or g13486 ( n13392 , n26519 , n3175 );
    or g13487 ( n15596 , n8493 , n16099 );
    xor g13488 ( n26433 , n8029 , n11204 );
    not g13489 ( n21159 , n7187 );
    xnor g13490 ( n14560 , n25884 , n9689 );
    or g13491 ( n24243 , n25466 , n21582 );
    and g13492 ( n8184 , n30136 , n13702 );
    or g13493 ( n13662 , n25789 , n700 );
    and g13494 ( n1023 , n28052 , n18588 );
    or g13495 ( n17186 , n26271 , n23618 );
    xnor g13496 ( n28624 , n6846 , n27112 );
    and g13497 ( n9843 , n2551 , n534 );
    xnor g13498 ( n23650 , n10559 , n13073 );
    xnor g13499 ( n20939 , n3410 , n21508 );
    or g13500 ( n9471 , n28445 , n8592 );
    and g13501 ( n12547 , n210 , n18661 );
    not g13502 ( n31228 , n28164 );
    not g13503 ( n9827 , n26500 );
    and g13504 ( n27122 , n9636 , n13514 );
    and g13505 ( n13789 , n4028 , n4103 );
    and g13506 ( n4415 , n22196 , n22394 );
    not g13507 ( n3280 , n31415 );
    or g13508 ( n4685 , n11837 , n10841 );
    xnor g13509 ( n28334 , n30242 , n15360 );
    xnor g13510 ( n23937 , n24784 , n26052 );
    and g13511 ( n4327 , n29488 , n22589 );
    not g13512 ( n22383 , n29380 );
    not g13513 ( n2154 , n17574 );
    and g13514 ( n15518 , n28519 , n24842 );
    not g13515 ( n1857 , n18804 );
    xnor g13516 ( n1131 , n1134 , n15922 );
    not g13517 ( n16106 , n25447 );
    and g13518 ( n24059 , n20163 , n3209 );
    nor g13519 ( n16600 , n18516 , n24402 );
    xnor g13520 ( n28564 , n13788 , n28311 );
    or g13521 ( n16504 , n8713 , n21243 );
    or g13522 ( n19075 , n30295 , n2233 );
    xor g13523 ( n25989 , n16863 , n30035 );
    not g13524 ( n31479 , n14962 );
    and g13525 ( n28798 , n20363 , n9100 );
    and g13526 ( n16926 , n8899 , n12424 );
    and g13527 ( n14552 , n16271 , n12784 );
    not g13528 ( n31653 , n26239 );
    not g13529 ( n4875 , n6295 );
    not g13530 ( n25821 , n22776 );
    or g13531 ( n1671 , n14255 , n29118 );
    or g13532 ( n5754 , n15825 , n9847 );
    nor g13533 ( n12612 , n17572 , n1614 );
    xnor g13534 ( n22257 , n7628 , n14243 );
    xnor g13535 ( n1088 , n20691 , n9626 );
    xnor g13536 ( n21133 , n3519 , n25276 );
    nor g13537 ( n80 , n12035 , n6775 );
    or g13538 ( n22580 , n28689 , n11422 );
    nor g13539 ( n4748 , n27233 , n29228 );
    nor g13540 ( n3889 , n419 , n16753 );
    or g13541 ( n5824 , n25516 , n4323 );
    or g13542 ( n20138 , n13629 , n29402 );
    nor g13543 ( n19665 , n28006 , n28449 );
    or g13544 ( n2935 , n25613 , n20028 );
    or g13545 ( n20401 , n29132 , n4122 );
    xnor g13546 ( n10741 , n20484 , n7776 );
    xnor g13547 ( n30838 , n9399 , n23411 );
    and g13548 ( n17372 , n23368 , n17368 );
    xnor g13549 ( n5967 , n24457 , n22408 );
    or g13550 ( n16682 , n1419 , n15437 );
    or g13551 ( n3170 , n26961 , n31668 );
    and g13552 ( n6860 , n28421 , n4485 );
    xnor g13553 ( n9805 , n23287 , n6325 );
    xnor g13554 ( n2313 , n13491 , n6460 );
    xnor g13555 ( n24544 , n9008 , n5251 );
    not g13556 ( n31309 , n15221 );
    and g13557 ( n14017 , n27319 , n27260 );
    or g13558 ( n8749 , n14226 , n15071 );
    or g13559 ( n11570 , n31027 , n29827 );
    not g13560 ( n11171 , n31591 );
    not g13561 ( n17693 , n7947 );
    not g13562 ( n19059 , n24696 );
    xnor g13563 ( n855 , n23325 , n25370 );
    or g13564 ( n14662 , n4769 , n5433 );
    and g13565 ( n8452 , n17546 , n12524 );
    xnor g13566 ( n28932 , n29513 , n18211 );
    not g13567 ( n9525 , n3095 );
    not g13568 ( n23277 , n20764 );
    or g13569 ( n25316 , n14572 , n16286 );
    not g13570 ( n19462 , n10731 );
    nor g13571 ( n28223 , n2924 , n26852 );
    not g13572 ( n8940 , n10913 );
    not g13573 ( n11226 , n27077 );
    and g13574 ( n28740 , n15445 , n19234 );
    or g13575 ( n5372 , n20529 , n26287 );
    xnor g13576 ( n6526 , n17273 , n27705 );
    xnor g13577 ( n27564 , n10984 , n30083 );
    xnor g13578 ( n6731 , n9022 , n21639 );
    or g13579 ( n27103 , n14421 , n15785 );
    and g13580 ( n21499 , n16749 , n26472 );
    and g13581 ( n24845 , n27332 , n31526 );
    and g13582 ( n25355 , n25729 , n11621 );
    or g13583 ( n32011 , n14992 , n742 );
    xnor g13584 ( n5833 , n7702 , n9633 );
    xor g13585 ( n10898 , n28407 , n17044 );
    xnor g13586 ( n31751 , n14286 , n28150 );
    xnor g13587 ( n31030 , n20883 , n27131 );
    or g13588 ( n17573 , n10061 , n19547 );
    xnor g13589 ( n6934 , n714 , n22728 );
    not g13590 ( n1002 , n30705 );
    not g13591 ( n3043 , n12803 );
    or g13592 ( n18049 , n1430 , n2014 );
    or g13593 ( n266 , n4716 , n17034 );
    xnor g13594 ( n29365 , n21180 , n1995 );
    not g13595 ( n7722 , n9467 );
    or g13596 ( n29251 , n23040 , n27936 );
    xnor g13597 ( n15143 , n30327 , n19630 );
    xnor g13598 ( n592 , n28807 , n8360 );
    xnor g13599 ( n16686 , n28158 , n23023 );
    or g13600 ( n23120 , n24333 , n23751 );
    not g13601 ( n12407 , n29923 );
    nor g13602 ( n13134 , n20390 , n20322 );
    xnor g13603 ( n23377 , n12280 , n11498 );
    not g13604 ( n6983 , n25793 );
    or g13605 ( n4365 , n28083 , n6314 );
    not g13606 ( n11764 , n9943 );
    xnor g13607 ( n4739 , n21729 , n8108 );
    xnor g13608 ( n4377 , n25182 , n27284 );
    and g13609 ( n24070 , n4954 , n15349 );
    xnor g13610 ( n5592 , n20278 , n21458 );
    not g13611 ( n21938 , n26568 );
    not g13612 ( n23786 , n23306 );
    xnor g13613 ( n5673 , n25937 , n1397 );
    or g13614 ( n9245 , n31381 , n15921 );
    or g13615 ( n18719 , n671 , n11514 );
    nor g13616 ( n26896 , n5022 , n28829 );
    nor g13617 ( n25349 , n8088 , n6281 );
    not g13618 ( n31916 , n9670 );
    nor g13619 ( n2797 , n22549 , n6896 );
    not g13620 ( n5378 , n22267 );
    xnor g13621 ( n21448 , n10034 , n28081 );
    or g13622 ( n2215 , n7514 , n26029 );
    not g13623 ( n25257 , n21307 );
    not g13624 ( n12758 , n3763 );
    or g13625 ( n1732 , n24221 , n6947 );
    not g13626 ( n7214 , n18825 );
    xnor g13627 ( n26999 , n22665 , n20815 );
    not g13628 ( n31091 , n30769 );
    and g13629 ( n25996 , n28500 , n256 );
    or g13630 ( n14642 , n2149 , n3308 );
    xnor g13631 ( n29242 , n9469 , n25291 );
    xnor g13632 ( n16389 , n21020 , n14252 );
    xnor g13633 ( n29843 , n20604 , n6525 );
    not g13634 ( n31973 , n3653 );
    not g13635 ( n22399 , n3163 );
    and g13636 ( n22611 , n10271 , n31696 );
    not g13637 ( n12986 , n752 );
    and g13638 ( n30302 , n28454 , n5002 );
    and g13639 ( n16802 , n11442 , n11570 );
    not g13640 ( n2473 , n15640 );
    not g13641 ( n4618 , n5388 );
    not g13642 ( n4730 , n9744 );
    or g13643 ( n10789 , n25572 , n3353 );
    nor g13644 ( n29033 , n3076 , n15568 );
    not g13645 ( n23285 , n20714 );
    and g13646 ( n29789 , n3129 , n30075 );
    not g13647 ( n22489 , n6306 );
    xnor g13648 ( n31757 , n2738 , n8402 );
    or g13649 ( n4025 , n7032 , n13946 );
    xnor g13650 ( n29972 , n23956 , n5511 );
    or g13651 ( n2002 , n2955 , n24307 );
    not g13652 ( n16111 , n1214 );
    xnor g13653 ( n9731 , n21636 , n19292 );
    or g13654 ( n24491 , n23138 , n29747 );
    and g13655 ( n7440 , n18006 , n21193 );
    xnor g13656 ( n19205 , n30524 , n24089 );
    not g13657 ( n12680 , n27706 );
    xnor g13658 ( n7278 , n7353 , n31283 );
    xor g13659 ( n10443 , n1555 , n23342 );
    not g13660 ( n31119 , n23047 );
    not g13661 ( n4176 , n17112 );
    and g13662 ( n7661 , n26626 , n2112 );
    or g13663 ( n9098 , n21929 , n23075 );
    or g13664 ( n2449 , n4563 , n30355 );
    not g13665 ( n28092 , n31347 );
    not g13666 ( n937 , n12668 );
    or g13667 ( n4682 , n19763 , n24054 );
    not g13668 ( n8725 , n29779 );
    and g13669 ( n6556 , n24495 , n9043 );
    xnor g13670 ( n10352 , n29935 , n8236 );
    and g13671 ( n14551 , n6548 , n14279 );
    or g13672 ( n4126 , n13866 , n12033 );
    or g13673 ( n13009 , n30014 , n2775 );
    xnor g13674 ( n7735 , n10338 , n22874 );
    and g13675 ( n27719 , n23279 , n20538 );
    not g13676 ( n10239 , n8875 );
    or g13677 ( n2030 , n26213 , n23671 );
    xnor g13678 ( n14806 , n2860 , n13611 );
    or g13679 ( n22833 , n10070 , n27902 );
    and g13680 ( n19468 , n8048 , n28125 );
    or g13681 ( n3027 , n6719 , n19457 );
    or g13682 ( n12698 , n26194 , n11397 );
    and g13683 ( n10666 , n16752 , n6631 );
    not g13684 ( n24696 , n28183 );
    not g13685 ( n4608 , n25089 );
    or g13686 ( n11568 , n3166 , n17784 );
    and g13687 ( n7006 , n7163 , n30838 );
    not g13688 ( n16409 , n5960 );
    not g13689 ( n30345 , n6695 );
    not g13690 ( n19184 , n31677 );
    not g13691 ( n16968 , n22734 );
    not g13692 ( n24873 , n12940 );
    and g13693 ( n26949 , n11113 , n9253 );
    not g13694 ( n29060 , n13410 );
    and g13695 ( n5160 , n27698 , n18826 );
    not g13696 ( n17761 , n20106 );
    nor g13697 ( n14001 , n10873 , n7557 );
    and g13698 ( n30447 , n30920 , n5308 );
    or g13699 ( n23737 , n7130 , n31004 );
    or g13700 ( n13456 , n23449 , n13854 );
    not g13701 ( n23153 , n13157 );
    nor g13702 ( n18347 , n4712 , n27696 );
    and g13703 ( n30027 , n23895 , n7554 );
    not g13704 ( n21621 , n58 );
    or g13705 ( n18006 , n12323 , n6710 );
    xnor g13706 ( n14663 , n24039 , n29153 );
    or g13707 ( n10663 , n8381 , n11021 );
    xnor g13708 ( n21865 , n5386 , n793 );
    not g13709 ( n29715 , n5628 );
    not g13710 ( n6858 , n13509 );
    or g13711 ( n876 , n16544 , n2667 );
    xor g13712 ( n16759 , n26358 , n27507 );
    not g13713 ( n19084 , n7381 );
    or g13714 ( n20133 , n19835 , n15457 );
    nor g13715 ( n25881 , n23638 , n29960 );
    and g13716 ( n13489 , n9226 , n2355 );
    or g13717 ( n15018 , n22253 , n31523 );
    or g13718 ( n570 , n14319 , n482 );
    not g13719 ( n8151 , n6424 );
    or g13720 ( n16801 , n8092 , n9171 );
    or g13721 ( n16107 , n8705 , n29918 );
    or g13722 ( n23186 , n30632 , n22657 );
    or g13723 ( n13071 , n3821 , n14689 );
    not g13724 ( n18057 , n1415 );
    xnor g13725 ( n7432 , n6795 , n29234 );
    or g13726 ( n23194 , n13038 , n30930 );
    xnor g13727 ( n4493 , n4494 , n30813 );
    not g13728 ( n19114 , n19322 );
    or g13729 ( n27874 , n1030 , n17062 );
    xnor g13730 ( n28320 , n30217 , n4587 );
    not g13731 ( n15491 , n23306 );
    and g13732 ( n21751 , n23661 , n27909 );
    and g13733 ( n5927 , n13658 , n26710 );
    not g13734 ( n29116 , n23536 );
    xnor g13735 ( n26785 , n27130 , n6949 );
    nor g13736 ( n489 , n6566 , n6070 );
    or g13737 ( n17361 , n20438 , n2813 );
    or g13738 ( n25255 , n15312 , n2886 );
    not g13739 ( n395 , n17454 );
    and g13740 ( n27288 , n19499 , n28586 );
    and g13741 ( n13651 , n14881 , n13969 );
    xnor g13742 ( n17591 , n10393 , n21597 );
    or g13743 ( n28224 , n30377 , n11681 );
    not g13744 ( n11540 , n5744 );
    xnor g13745 ( n31002 , n24719 , n28822 );
    xnor g13746 ( n16314 , n21022 , n2676 );
    and g13747 ( n3442 , n160 , n30008 );
    or g13748 ( n877 , n31018 , n4200 );
    not g13749 ( n5917 , n3682 );
    not g13750 ( n30623 , n23635 );
    xnor g13751 ( n796 , n18351 , n5570 );
    not g13752 ( n24294 , n100 );
    and g13753 ( n20188 , n2696 , n30081 );
    nor g13754 ( n5320 , n9652 , n21833 );
    and g13755 ( n25812 , n3379 , n11739 );
    xor g13756 ( n5941 , n11207 , n20194 );
    or g13757 ( n16440 , n18229 , n7859 );
    xnor g13758 ( n13280 , n13827 , n6143 );
    and g13759 ( n4250 , n19971 , n26272 );
    and g13760 ( n8288 , n3120 , n12583 );
    nor g13761 ( n23754 , n22398 , n2657 );
    or g13762 ( n5347 , n15013 , n27641 );
    not g13763 ( n9078 , n31455 );
    nor g13764 ( n1862 , n23735 , n16660 );
    xnor g13765 ( n4832 , n30388 , n897 );
    not g13766 ( n3342 , n17823 );
    xnor g13767 ( n22490 , n19289 , n28659 );
    or g13768 ( n11876 , n19066 , n19516 );
    and g13769 ( n27105 , n6029 , n8656 );
    xnor g13770 ( n6564 , n29488 , n2913 );
    or g13771 ( n22303 , n8279 , n12350 );
    not g13772 ( n19489 , n10443 );
    xnor g13773 ( n20679 , n5120 , n7884 );
    not g13774 ( n15151 , n19852 );
    or g13775 ( n10192 , n22532 , n24027 );
    or g13776 ( n19725 , n22451 , n28222 );
    xnor g13777 ( n26771 , n31849 , n29380 );
    not g13778 ( n31359 , n6766 );
    xnor g13779 ( n6274 , n27080 , n19358 );
    or g13780 ( n13490 , n31320 , n19894 );
    xor g13781 ( n30798 , n26567 , n23208 );
    xnor g13782 ( n30250 , n15575 , n17665 );
    xnor g13783 ( n10289 , n11432 , n31079 );
    or g13784 ( n4905 , n14752 , n15225 );
    xnor g13785 ( n8428 , n12400 , n513 );
    not g13786 ( n23497 , n29961 );
    not g13787 ( n29714 , n2177 );
    or g13788 ( n20670 , n23418 , n27859 );
    and g13789 ( n27765 , n14378 , n21489 );
    xnor g13790 ( n24591 , n30443 , n31927 );
    xnor g13791 ( n20249 , n26454 , n138 );
    xnor g13792 ( n3006 , n8063 , n30534 );
    xnor g13793 ( n11194 , n27175 , n26763 );
    not g13794 ( n28607 , n20964 );
    not g13795 ( n12448 , n22754 );
    not g13796 ( n27570 , n20505 );
    not g13797 ( n15640 , n23029 );
    and g13798 ( n29805 , n11447 , n1141 );
    and g13799 ( n23880 , n14632 , n25676 );
    not g13800 ( n25835 , n11730 );
    or g13801 ( n25990 , n23062 , n28567 );
    nor g13802 ( n17101 , n8166 , n6983 );
    nor g13803 ( n19058 , n23608 , n5443 );
    xnor g13804 ( n20096 , n14690 , n10269 );
    and g13805 ( n13107 , n9722 , n27458 );
    or g13806 ( n13465 , n16558 , n26373 );
    not g13807 ( n10799 , n28837 );
    nor g13808 ( n9861 , n16148 , n17632 );
    not g13809 ( n16392 , n2032 );
    and g13810 ( n12945 , n6894 , n371 );
    not g13811 ( n5964 , n19035 );
    or g13812 ( n2501 , n27147 , n27763 );
    not g13813 ( n8736 , n12325 );
    nor g13814 ( n20876 , n13751 , n16625 );
    xor g13815 ( n16778 , n10604 , n21490 );
    not g13816 ( n3735 , n12056 );
    xnor g13817 ( n17257 , n16073 , n29631 );
    xnor g13818 ( n18360 , n8141 , n24569 );
    not g13819 ( n13744 , n6280 );
    or g13820 ( n28208 , n13496 , n17635 );
    xnor g13821 ( n29360 , n19060 , n14208 );
    or g13822 ( n8773 , n28862 , n9052 );
    not g13823 ( n16574 , n27022 );
    or g13824 ( n22152 , n26823 , n23343 );
    xnor g13825 ( n28533 , n2586 , n25579 );
    xnor g13826 ( n15340 , n575 , n25261 );
    not g13827 ( n16914 , n12207 );
    not g13828 ( n22591 , n22546 );
    or g13829 ( n14301 , n10388 , n25392 );
    or g13830 ( n31734 , n862 , n22605 );
    not g13831 ( n13086 , n25569 );
    xnor g13832 ( n21106 , n23442 , n2090 );
    not g13833 ( n19324 , n5985 );
    or g13834 ( n16566 , n20637 , n24645 );
    xnor g13835 ( n24664 , n260 , n7296 );
    or g13836 ( n7911 , n6997 , n27554 );
    nor g13837 ( n30152 , n14121 , n7009 );
    or g13838 ( n23210 , n30663 , n28359 );
    not g13839 ( n10794 , n13492 );
    xnor g13840 ( n22361 , n1151 , n14627 );
    and g13841 ( n27558 , n16277 , n6256 );
    xnor g13842 ( n17695 , n14347 , n10741 );
    and g13843 ( n2733 , n7916 , n7300 );
    not g13844 ( n2112 , n15 );
    xnor g13845 ( n17993 , n16284 , n10696 );
    xnor g13846 ( n1254 , n28084 , n2825 );
    xnor g13847 ( n10014 , n25722 , n27777 );
    xnor g13848 ( n31365 , n17758 , n7655 );
    xnor g13849 ( n3524 , n24427 , n6950 );
    nor g13850 ( n4846 , n22514 , n9473 );
    not g13851 ( n26286 , n14005 );
    nor g13852 ( n20324 , n4662 , n17514 );
    nor g13853 ( n15686 , n26888 , n1179 );
    nor g13854 ( n2214 , n17032 , n28315 );
    xnor g13855 ( n2467 , n26081 , n21885 );
    and g13856 ( n21406 , n18171 , n16150 );
    xnor g13857 ( n30566 , n12414 , n1858 );
    xnor g13858 ( n9234 , n4635 , n2316 );
    nor g13859 ( n18584 , n8898 , n22141 );
    xnor g13860 ( n17058 , n15775 , n14980 );
    and g13861 ( n14543 , n24046 , n13419 );
    and g13862 ( n15955 , n28788 , n26174 );
    xnor g13863 ( n10456 , n29990 , n14190 );
    xnor g13864 ( n11716 , n29518 , n8344 );
    and g13865 ( n23359 , n390 , n14597 );
    or g13866 ( n11320 , n26367 , n29135 );
    or g13867 ( n4265 , n5594 , n8999 );
    and g13868 ( n3908 , n4603 , n1235 );
    and g13869 ( n22506 , n29621 , n2349 );
    not g13870 ( n16602 , n10013 );
    or g13871 ( n26981 , n20041 , n2311 );
    xnor g13872 ( n24338 , n2307 , n1246 );
    not g13873 ( n986 , n31287 );
    nor g13874 ( n19603 , n4844 , n19538 );
    and g13875 ( n4752 , n31760 , n21456 );
    xnor g13876 ( n28835 , n12771 , n5149 );
    and g13877 ( n699 , n5482 , n16251 );
    xnor g13878 ( n28124 , n14442 , n20716 );
    not g13879 ( n14547 , n10153 );
    xnor g13880 ( n8336 , n3098 , n89 );
    not g13881 ( n9087 , n31878 );
    or g13882 ( n30986 , n15734 , n23693 );
    xnor g13883 ( n11614 , n18481 , n3815 );
    and g13884 ( n6587 , n25015 , n28122 );
    or g13885 ( n1741 , n19027 , n23393 );
    or g13886 ( n24030 , n17327 , n26967 );
    not g13887 ( n21631 , n1606 );
    and g13888 ( n10840 , n20602 , n20548 );
    and g13889 ( n4360 , n7650 , n198 );
    xnor g13890 ( n111 , n25092 , n31556 );
    and g13891 ( n53 , n6156 , n5096 );
    not g13892 ( n3864 , n16250 );
    not g13893 ( n6152 , n29301 );
    xnor g13894 ( n20359 , n28769 , n11457 );
    nor g13895 ( n1939 , n7355 , n302 );
    not g13896 ( n25613 , n17653 );
    or g13897 ( n8992 , n6236 , n5065 );
    or g13898 ( n22511 , n15796 , n12019 );
    or g13899 ( n23553 , n2980 , n27428 );
    or g13900 ( n15327 , n24229 , n1363 );
    or g13901 ( n11364 , n15381 , n26744 );
    or g13902 ( n17066 , n14106 , n20748 );
    and g13903 ( n14768 , n24878 , n12947 );
    not g13904 ( n24698 , n8574 );
    and g13905 ( n5549 , n3448 , n20314 );
    not g13906 ( n15275 , n6437 );
    and g13907 ( n2201 , n1655 , n15811 );
    not g13908 ( n13684 , n31306 );
    or g13909 ( n12531 , n24195 , n23253 );
    not g13910 ( n14405 , n7336 );
    not g13911 ( n7524 , n9401 );
    or g13912 ( n31668 , n27034 , n29059 );
    nor g13913 ( n3750 , n17109 , n30632 );
    and g13914 ( n14502 , n7072 , n10248 );
    nor g13915 ( n18138 , n23043 , n10931 );
    nor g13916 ( n2765 , n18067 , n30262 );
    xnor g13917 ( n6639 , n11596 , n5916 );
    or g13918 ( n15063 , n6046 , n4299 );
    and g13919 ( n21414 , n13803 , n27082 );
    xnor g13920 ( n5144 , n28417 , n9691 );
    or g13921 ( n23792 , n3385 , n8966 );
    xnor g13922 ( n13854 , n14179 , n20384 );
    and g13923 ( n26330 , n6097 , n19708 );
    xnor g13924 ( n15418 , n22917 , n3080 );
    not g13925 ( n16284 , n15472 );
    or g13926 ( n25977 , n16238 , n12031 );
    not g13927 ( n28768 , n15906 );
    xnor g13928 ( n10836 , n12072 , n18534 );
    nor g13929 ( n11727 , n17130 , n27172 );
    xnor g13930 ( n29684 , n25991 , n19217 );
    not g13931 ( n20452 , n18371 );
    not g13932 ( n12022 , n10542 );
    nor g13933 ( n24064 , n29397 , n11640 );
    not g13934 ( n15530 , n16741 );
    and g13935 ( n27314 , n21471 , n15058 );
    not g13936 ( n4916 , n19443 );
    or g13937 ( n29783 , n393 , n8826 );
    xnor g13938 ( n9368 , n24970 , n11313 );
    and g13939 ( n26688 , n20818 , n24604 );
    xnor g13940 ( n2502 , n3307 , n12514 );
    or g13941 ( n28056 , n2444 , n24916 );
    not g13942 ( n8582 , n31387 );
    not g13943 ( n2720 , n26966 );
    not g13944 ( n28755 , n27106 );
    not g13945 ( n11234 , n26268 );
    or g13946 ( n30284 , n9372 , n15426 );
    and g13947 ( n29383 , n4406 , n14353 );
    nor g13948 ( n25572 , n29818 , n4956 );
    or g13949 ( n18796 , n20070 , n9240 );
    not g13950 ( n21669 , n12178 );
    not g13951 ( n15431 , n25276 );
    not g13952 ( n14952 , n22371 );
    not g13953 ( n19679 , n30427 );
    xnor g13954 ( n17328 , n12958 , n24607 );
    xnor g13955 ( n14131 , n18689 , n31512 );
    nor g13956 ( n30309 , n3782 , n13510 );
    not g13957 ( n7798 , n26580 );
    not g13958 ( n11595 , n1521 );
    xnor g13959 ( n20914 , n11474 , n18116 );
    not g13960 ( n16586 , n22505 );
    xnor g13961 ( n11915 , n20495 , n30525 );
    or g13962 ( n16305 , n6601 , n1313 );
    nor g13963 ( n27273 , n16412 , n31652 );
    xnor g13964 ( n18755 , n20573 , n8360 );
    or g13965 ( n759 , n30651 , n1794 );
    not g13966 ( n3046 , n21282 );
    and g13967 ( n11106 , n11530 , n15561 );
    and g13968 ( n8199 , n23904 , n8755 );
    or g13969 ( n9140 , n17177 , n21446 );
    xnor g13970 ( n18108 , n26117 , n2939 );
    and g13971 ( n14862 , n16323 , n28358 );
    not g13972 ( n19704 , n6703 );
    and g13973 ( n15704 , n15294 , n20239 );
    xnor g13974 ( n13028 , n21394 , n30865 );
    not g13975 ( n20066 , n1880 );
    or g13976 ( n12915 , n10779 , n13893 );
    nor g13977 ( n26821 , n10772 , n9538 );
    and g13978 ( n30899 , n20459 , n30242 );
    nor g13979 ( n24044 , n23114 , n17795 );
    or g13980 ( n3802 , n6181 , n30988 );
    and g13981 ( n15641 , n27519 , n31670 );
    xor g13982 ( n12325 , n3992 , n10139 );
    xnor g13983 ( n1126 , n18127 , n13846 );
    nor g13984 ( n145 , n15140 , n30327 );
    and g13985 ( n18560 , n9125 , n10725 );
    and g13986 ( n12416 , n8205 , n10513 );
    not g13987 ( n4968 , n6707 );
    nor g13988 ( n1217 , n11065 , n28979 );
    and g13989 ( n15002 , n26443 , n516 );
    or g13990 ( n10892 , n31876 , n21799 );
    xnor g13991 ( n23309 , n28907 , n20158 );
    and g13992 ( n26865 , n31705 , n29082 );
    not g13993 ( n15142 , n30908 );
    or g13994 ( n31457 , n3339 , n29225 );
    not g13995 ( n8423 , n18645 );
    not g13996 ( n28245 , n16558 );
    not g13997 ( n28709 , n17265 );
    or g13998 ( n13409 , n398 , n15419 );
    and g13999 ( n22347 , n27113 , n13006 );
    not g14000 ( n10146 , n8256 );
    and g14001 ( n4426 , n25350 , n14533 );
    and g14002 ( n421 , n8124 , n7701 );
    or g14003 ( n15817 , n5837 , n29716 );
    xnor g14004 ( n779 , n8042 , n29249 );
    xor g14005 ( n31996 , n15828 , n20304 );
    or g14006 ( n11380 , n18566 , n24207 );
    and g14007 ( n20323 , n28312 , n24511 );
    not g14008 ( n6024 , n10236 );
    xnor g14009 ( n16677 , n23051 , n25636 );
    not g14010 ( n4172 , n19067 );
    xnor g14011 ( n11971 , n14477 , n19956 );
    xnor g14012 ( n25783 , n18389 , n1039 );
    or g14013 ( n12393 , n2792 , n17306 );
    xnor g14014 ( n22642 , n13132 , n8009 );
    not g14015 ( n14604 , n3641 );
    or g14016 ( n30877 , n29821 , n29034 );
    nor g14017 ( n14393 , n25319 , n7446 );
    xnor g14018 ( n11782 , n5461 , n17687 );
    or g14019 ( n16553 , n25948 , n130 );
    and g14020 ( n12058 , n28064 , n17980 );
    xnor g14021 ( n7384 , n24348 , n28739 );
    or g14022 ( n20054 , n26822 , n22983 );
    or g14023 ( n4185 , n4554 , n11204 );
    not g14024 ( n24709 , n3846 );
    and g14025 ( n4654 , n14042 , n8112 );
    nor g14026 ( n26691 , n19132 , n31259 );
    or g14027 ( n30926 , n14062 , n3116 );
    not g14028 ( n21710 , n25756 );
    xnor g14029 ( n20771 , n15247 , n26604 );
    xnor g14030 ( n1770 , n28235 , n10623 );
    and g14031 ( n11865 , n17047 , n25736 );
    or g14032 ( n28696 , n23876 , n24287 );
    not g14033 ( n15253 , n7896 );
    xnor g14034 ( n10335 , n29750 , n27767 );
    not g14035 ( n4050 , n5853 );
    xnor g14036 ( n14430 , n27941 , n14658 );
    or g14037 ( n27231 , n27681 , n26806 );
    nor g14038 ( n16435 , n13939 , n12519 );
    or g14039 ( n1315 , n3810 , n11180 );
    not g14040 ( n925 , n12188 );
    xnor g14041 ( n2758 , n25276 , n4844 );
    not g14042 ( n15328 , n13839 );
    not g14043 ( n10411 , n21767 );
    or g14044 ( n2327 , n17794 , n31335 );
    not g14045 ( n4476 , n30741 );
    or g14046 ( n20635 , n9915 , n17432 );
    xnor g14047 ( n21389 , n22054 , n523 );
    xnor g14048 ( n22747 , n53 , n22455 );
    xnor g14049 ( n12595 , n2542 , n9486 );
    not g14050 ( n22042 , n16943 );
    nor g14051 ( n30972 , n18391 , n27233 );
    nor g14052 ( n15555 , n29060 , n4786 );
    and g14053 ( n5777 , n30993 , n5713 );
    and g14054 ( n656 , n26334 , n19782 );
    xnor g14055 ( n14272 , n6666 , n26414 );
    or g14056 ( n24460 , n22360 , n16121 );
    not g14057 ( n28630 , n15610 );
    xnor g14058 ( n3621 , n2213 , n2686 );
    or g14059 ( n24872 , n27868 , n19044 );
    xnor g14060 ( n2054 , n22648 , n12329 );
    xnor g14061 ( n14929 , n621 , n16516 );
    or g14062 ( n27544 , n24035 , n30763 );
    or g14063 ( n31656 , n27741 , n12569 );
    not g14064 ( n1273 , n21261 );
    nor g14065 ( n9844 , n16481 , n16651 );
    xnor g14066 ( n9480 , n10257 , n24315 );
    xnor g14067 ( n24965 , n4893 , n28583 );
    xnor g14068 ( n29303 , n12025 , n2386 );
    and g14069 ( n17592 , n3639 , n25699 );
    or g14070 ( n25719 , n17019 , n30853 );
    not g14071 ( n7682 , n10289 );
    or g14072 ( n18231 , n14937 , n12775 );
    or g14073 ( n20016 , n9653 , n18040 );
    not g14074 ( n7757 , n7760 );
    and g14075 ( n732 , n28568 , n8590 );
    xnor g14076 ( n9729 , n30332 , n3417 );
    or g14077 ( n13929 , n10474 , n27135 );
    xnor g14078 ( n10113 , n9116 , n12030 );
    xnor g14079 ( n4247 , n11538 , n17705 );
    nor g14080 ( n29138 , n30732 , n25761 );
    or g14081 ( n26757 , n916 , n30698 );
    not g14082 ( n25031 , n17006 );
    xor g14083 ( n3854 , n27168 , n12514 );
    and g14084 ( n29907 , n22971 , n2097 );
    nor g14085 ( n19838 , n3106 , n9412 );
    xor g14086 ( n19721 , n8287 , n17559 );
    not g14087 ( n27997 , n4739 );
    not g14088 ( n29400 , n8714 );
    not g14089 ( n23010 , n12388 );
    and g14090 ( n11022 , n22317 , n27923 );
    and g14091 ( n16133 , n5157 , n538 );
    not g14092 ( n7154 , n579 );
    and g14093 ( n11563 , n20026 , n16535 );
    xor g14094 ( n15492 , n3060 , n7095 );
    xnor g14095 ( n15810 , n3954 , n28685 );
    not g14096 ( n11514 , n1020 );
    or g14097 ( n26480 , n30832 , n14775 );
    and g14098 ( n19431 , n2801 , n24837 );
    and g14099 ( n9297 , n17843 , n15758 );
    xnor g14100 ( n20082 , n31764 , n20577 );
    and g14101 ( n17565 , n30774 , n16662 );
    or g14102 ( n21433 , n1935 , n5876 );
    xnor g14103 ( n5684 , n13534 , n3828 );
    xnor g14104 ( n22262 , n22181 , n4861 );
    not g14105 ( n13319 , n23844 );
    not g14106 ( n10228 , n20632 );
    nor g14107 ( n3893 , n21377 , n1485 );
    nor g14108 ( n1437 , n13463 , n23276 );
    xnor g14109 ( n18007 , n8119 , n31637 );
    nor g14110 ( n13366 , n24323 , n9905 );
    not g14111 ( n30244 , n27077 );
    xnor g14112 ( n1628 , n30769 , n11643 );
    xnor g14113 ( n9611 , n12452 , n31515 );
    xnor g14114 ( n11552 , n5761 , n10544 );
    or g14115 ( n25723 , n27026 , n358 );
    and g14116 ( n24936 , n21074 , n23961 );
    not g14117 ( n11836 , n18192 );
    xnor g14118 ( n2277 , n6070 , n23044 );
    and g14119 ( n21656 , n13618 , n166 );
    and g14120 ( n25548 , n29125 , n15557 );
    xnor g14121 ( n9092 , n664 , n9414 );
    not g14122 ( n16129 , n28597 );
    not g14123 ( n12440 , n1449 );
    xnor g14124 ( n431 , n5141 , n8780 );
    not g14125 ( n2213 , n12182 );
    or g14126 ( n24941 , n27064 , n8873 );
    xnor g14127 ( n26299 , n31509 , n13837 );
    or g14128 ( n18801 , n413 , n18567 );
    not g14129 ( n11663 , n8397 );
    not g14130 ( n21030 , n22917 );
    xnor g14131 ( n12049 , n1631 , n13644 );
    or g14132 ( n26978 , n2547 , n1109 );
    and g14133 ( n22680 , n25456 , n29251 );
    not g14134 ( n17317 , n19062 );
    and g14135 ( n15119 , n24381 , n9939 );
    not g14136 ( n28588 , n27127 );
    not g14137 ( n20110 , n15269 );
    xor g14138 ( n17398 , n12983 , n953 );
    not g14139 ( n17503 , n7907 );
    xnor g14140 ( n28431 , n10281 , n12960 );
    xnor g14141 ( n9062 , n27853 , n8898 );
    xnor g14142 ( n13135 , n13969 , n31355 );
    not g14143 ( n28139 , n26277 );
    not g14144 ( n9549 , n30936 );
    not g14145 ( n5566 , n10703 );
    nor g14146 ( n28921 , n5387 , n3639 );
    or g14147 ( n2917 , n23909 , n16954 );
    xnor g14148 ( n8792 , n25024 , n9478 );
    or g14149 ( n15503 , n19935 , n8403 );
    or g14150 ( n20201 , n22262 , n27996 );
    or g14151 ( n8648 , n674 , n4383 );
    or g14152 ( n30977 , n31431 , n30373 );
    xnor g14153 ( n31027 , n32017 , n29126 );
    or g14154 ( n3301 , n11362 , n20270 );
    or g14155 ( n27156 , n25747 , n17162 );
    or g14156 ( n6514 , n31636 , n18721 );
    not g14157 ( n18283 , n13451 );
    nor g14158 ( n9685 , n1176 , n21768 );
    nor g14159 ( n23362 , n16676 , n2779 );
    or g14160 ( n10903 , n680 , n2931 );
    not g14161 ( n20644 , n20181 );
    buf g14162 ( n11110 , n23716 );
    or g14163 ( n4387 , n14306 , n8038 );
    xnor g14164 ( n18933 , n24265 , n1531 );
    not g14165 ( n10368 , n29274 );
    xnor g14166 ( n9643 , n11431 , n20531 );
    and g14167 ( n24840 , n4036 , n30521 );
    xnor g14168 ( n14235 , n8756 , n23486 );
    and g14169 ( n10059 , n1240 , n18650 );
    nor g14170 ( n11505 , n18451 , n19556 );
    xnor g14171 ( n24660 , n27047 , n18823 );
    and g14172 ( n18961 , n16051 , n27557 );
    xnor g14173 ( n15986 , n18642 , n7698 );
    not g14174 ( n15604 , n25527 );
    or g14175 ( n26815 , n24327 , n2255 );
    not g14176 ( n3387 , n26610 );
    or g14177 ( n29455 , n18238 , n1181 );
    or g14178 ( n31341 , n31467 , n17990 );
    not g14179 ( n15055 , n7033 );
    or g14180 ( n31565 , n5617 , n29955 );
    or g14181 ( n16184 , n14351 , n24738 );
    or g14182 ( n14396 , n31293 , n16960 );
    not g14183 ( n17267 , n23496 );
    xnor g14184 ( n25826 , n30807 , n1946 );
    xnor g14185 ( n4239 , n6751 , n19701 );
    not g14186 ( n9500 , n6754 );
    xnor g14187 ( n21806 , n104 , n20952 );
    xnor g14188 ( n25380 , n7854 , n23189 );
    not g14189 ( n30587 , n10686 );
    or g14190 ( n22026 , n24695 , n10147 );
    and g14191 ( n18330 , n27115 , n2200 );
    xnor g14192 ( n7899 , n28532 , n13648 );
    or g14193 ( n15099 , n27546 , n1230 );
    not g14194 ( n30822 , n19572 );
    and g14195 ( n6617 , n19307 , n7443 );
    xnor g14196 ( n17472 , n31498 , n24066 );
    and g14197 ( n27640 , n1136 , n30109 );
    or g14198 ( n22999 , n5131 , n25808 );
    not g14199 ( n17448 , n15891 );
    and g14200 ( n1984 , n13874 , n11145 );
    or g14201 ( n23244 , n21902 , n20888 );
    or g14202 ( n19342 , n26665 , n18068 );
    not g14203 ( n3406 , n31026 );
    nor g14204 ( n31122 , n22399 , n20922 );
    nor g14205 ( n14659 , n9529 , n2800 );
    or g14206 ( n1300 , n19497 , n5463 );
    not g14207 ( n15495 , n24939 );
    nor g14208 ( n895 , n24512 , n2872 );
    not g14209 ( n17183 , n9820 );
    or g14210 ( n29205 , n17798 , n26378 );
    not g14211 ( n4004 , n24137 );
    or g14212 ( n19441 , n19023 , n8399 );
    nor g14213 ( n8535 , n22233 , n25760 );
    xnor g14214 ( n9215 , n13908 , n10841 );
    not g14215 ( n22647 , n11414 );
    or g14216 ( n17787 , n8764 , n12851 );
    xnor g14217 ( n28227 , n10371 , n1562 );
    nor g14218 ( n6099 , n5036 , n26026 );
    not g14219 ( n26459 , n5679 );
    not g14220 ( n26116 , n27595 );
    not g14221 ( n858 , n21685 );
    buf g14222 ( n14376 , n7064 );
    nor g14223 ( n31525 , n27896 , n11610 );
    not g14224 ( n20468 , n22919 );
    not g14225 ( n25595 , n10959 );
    or g14226 ( n3250 , n22178 , n2323 );
    xnor g14227 ( n29467 , n2798 , n17499 );
    not g14228 ( n10712 , n10689 );
    or g14229 ( n30416 , n11720 , n17155 );
    xnor g14230 ( n28598 , n18695 , n16267 );
    not g14231 ( n12926 , n2070 );
    xnor g14232 ( n6852 , n13833 , n22512 );
    nor g14233 ( n5604 , n18234 , n31880 );
    not g14234 ( n29803 , n16956 );
    and g14235 ( n12471 , n97 , n21918 );
    or g14236 ( n8868 , n25130 , n6246 );
    or g14237 ( n31756 , n26374 , n25492 );
    nor g14238 ( n14728 , n12475 , n7431 );
    not g14239 ( n22906 , n2106 );
    or g14240 ( n822 , n15860 , n15310 );
    not g14241 ( n21803 , n27537 );
    not g14242 ( n4714 , n11944 );
    xnor g14243 ( n19105 , n9840 , n29190 );
    and g14244 ( n7507 , n15785 , n387 );
    or g14245 ( n26045 , n8682 , n24092 );
    or g14246 ( n10722 , n14114 , n7526 );
    xnor g14247 ( n29691 , n27212 , n14870 );
    or g14248 ( n22054 , n15497 , n16926 );
    not g14249 ( n11157 , n20803 );
    not g14250 ( n19814 , n5544 );
    xnor g14251 ( n16860 , n27136 , n14911 );
    and g14252 ( n3878 , n5245 , n13223 );
    xor g14253 ( n17165 , n18109 , n19785 );
    not g14254 ( n12993 , n19068 );
    or g14255 ( n31629 , n5570 , n24308 );
    or g14256 ( n9183 , n31476 , n9557 );
    not g14257 ( n423 , n11906 );
    nor g14258 ( n3896 , n17051 , n12277 );
    or g14259 ( n4975 , n26711 , n21002 );
    or g14260 ( n28714 , n6042 , n15675 );
    or g14261 ( n12395 , n6471 , n5017 );
    and g14262 ( n31496 , n19050 , n30607 );
    and g14263 ( n7724 , n15564 , n24756 );
    xnor g14264 ( n10889 , n8714 , n5873 );
    nor g14265 ( n30179 , n23101 , n21228 );
    and g14266 ( n7239 , n3823 , n15047 );
    and g14267 ( n8941 , n3873 , n10737 );
    and g14268 ( n21295 , n21771 , n17227 );
    xnor g14269 ( n26391 , n4552 , n2403 );
    not g14270 ( n6245 , n28766 );
    not g14271 ( n30546 , n1720 );
    and g14272 ( n5450 , n26104 , n29597 );
    or g14273 ( n3882 , n14274 , n3677 );
    xnor g14274 ( n22085 , n20739 , n24775 );
    xnor g14275 ( n865 , n577 , n31622 );
    not g14276 ( n30094 , n19407 );
    nor g14277 ( n4931 , n11494 , n28105 );
    nor g14278 ( n5954 , n1348 , n17927 );
    xnor g14279 ( n14864 , n11435 , n12141 );
    xnor g14280 ( n15059 , n26776 , n17932 );
    not g14281 ( n19492 , n31051 );
    xnor g14282 ( n5686 , n18925 , n22447 );
    xnor g14283 ( n14190 , n28929 , n25566 );
    or g14284 ( n8048 , n26643 , n2947 );
    and g14285 ( n29034 , n28265 , n24752 );
    not g14286 ( n29253 , n906 );
    xnor g14287 ( n9111 , n7434 , n30908 );
    or g14288 ( n21488 , n22944 , n31558 );
    or g14289 ( n9694 , n30700 , n8708 );
    and g14290 ( n18172 , n18341 , n31272 );
    and g14291 ( n4273 , n22596 , n12556 );
    or g14292 ( n30480 , n346 , n29842 );
    or g14293 ( n30715 , n30915 , n18468 );
    or g14294 ( n11862 , n6416 , n30238 );
    or g14295 ( n25229 , n11867 , n31483 );
    xnor g14296 ( n27742 , n10561 , n20412 );
    nor g14297 ( n16875 , n13935 , n4535 );
    or g14298 ( n15979 , n126 , n425 );
    and g14299 ( n30508 , n24472 , n30854 );
    and g14300 ( n11603 , n5931 , n3358 );
    and g14301 ( n28099 , n4184 , n16488 );
    not g14302 ( n25761 , n1688 );
    or g14303 ( n6920 , n15722 , n12863 );
    or g14304 ( n13986 , n4961 , n15786 );
    and g14305 ( n1621 , n1117 , n2400 );
    not g14306 ( n24196 , n14563 );
    or g14307 ( n15352 , n19217 , n24173 );
    or g14308 ( n22230 , n23240 , n21179 );
    xnor g14309 ( n12322 , n11355 , n624 );
    not g14310 ( n31419 , n24325 );
    not g14311 ( n5356 , n10231 );
    and g14312 ( n310 , n3263 , n27749 );
    not g14313 ( n23341 , n15252 );
    not g14314 ( n30349 , n11070 );
    nor g14315 ( n7027 , n16214 , n30739 );
    and g14316 ( n3155 , n17164 , n15172 );
    not g14317 ( n23332 , n11211 );
    xnor g14318 ( n22851 , n5895 , n28417 );
    or g14319 ( n17809 , n13640 , n23893 );
    or g14320 ( n30702 , n20234 , n6956 );
    and g14321 ( n2922 , n4392 , n25949 );
    xnor g14322 ( n11430 , n26974 , n16986 );
    and g14323 ( n28805 , n5139 , n7339 );
    xnor g14324 ( n29072 , n27513 , n17651 );
    or g14325 ( n1555 , n2248 , n24589 );
    or g14326 ( n29273 , n3152 , n21393 );
    nor g14327 ( n22562 , n2705 , n15892 );
    not g14328 ( n2684 , n483 );
    xnor g14329 ( n20039 , n2170 , n17919 );
    not g14330 ( n29539 , n11148 );
    or g14331 ( n5370 , n30068 , n26040 );
    or g14332 ( n5693 , n11236 , n4428 );
    nor g14333 ( n3690 , n30525 , n5711 );
    and g14334 ( n28581 , n25876 , n23194 );
    or g14335 ( n1460 , n6627 , n8679 );
    not g14336 ( n12195 , n16558 );
    and g14337 ( n16162 , n848 , n31317 );
    not g14338 ( n2982 , n23455 );
    nor g14339 ( n28687 , n22652 , n6361 );
    not g14340 ( n1302 , n20799 );
    nor g14341 ( n31475 , n14292 , n29890 );
    nor g14342 ( n21600 , n27491 , n7937 );
    not g14343 ( n551 , n18907 );
    and g14344 ( n6479 , n15350 , n29167 );
    not g14345 ( n24331 , n14520 );
    nor g14346 ( n964 , n20528 , n11106 );
    xnor g14347 ( n24769 , n5718 , n6909 );
    not g14348 ( n31755 , n21584 );
    xor g14349 ( n3276 , n21284 , n21497 );
    xnor g14350 ( n27359 , n25834 , n7993 );
    xnor g14351 ( n9984 , n14500 , n28932 );
    not g14352 ( n11765 , n7851 );
    xnor g14353 ( n17504 , n24465 , n24837 );
    xnor g14354 ( n12704 , n17936 , n20679 );
    and g14355 ( n17593 , n24180 , n22234 );
    xnor g14356 ( n18065 , n10170 , n31210 );
    or g14357 ( n14234 , n31498 , n19364 );
    or g14358 ( n11318 , n1417 , n4883 );
    and g14359 ( n24139 , n344 , n179 );
    or g14360 ( n18742 , n511 , n3092 );
    or g14361 ( n20542 , n3206 , n4544 );
    and g14362 ( n11900 , n26762 , n24894 );
    nor g14363 ( n24394 , n10851 , n21566 );
    and g14364 ( n16994 , n12994 , n26867 );
    xnor g14365 ( n26474 , n23852 , n14290 );
    or g14366 ( n9065 , n25703 , n24466 );
    not g14367 ( n31288 , n25242 );
    or g14368 ( n28706 , n1005 , n7460 );
    not g14369 ( n19041 , n23216 );
    and g14370 ( n24760 , n2839 , n22066 );
    or g14371 ( n25207 , n9736 , n2710 );
    and g14372 ( n26273 , n27479 , n15768 );
    xnor g14373 ( n28034 , n28568 , n11549 );
    not g14374 ( n4122 , n25976 );
    not g14375 ( n518 , n10827 );
    and g14376 ( n25289 , n18335 , n27282 );
    xnor g14377 ( n6610 , n24505 , n17394 );
    and g14378 ( n1168 , n21617 , n10782 );
    or g14379 ( n5572 , n18698 , n1693 );
    xnor g14380 ( n2056 , n6303 , n6727 );
    or g14381 ( n3437 , n17067 , n9713 );
    or g14382 ( n12164 , n27745 , n25932 );
    or g14383 ( n19685 , n14336 , n1288 );
    xnor g14384 ( n16071 , n20002 , n3720 );
    xnor g14385 ( n28901 , n16865 , n26264 );
    buf g14386 ( n2386 , n9317 );
    xnor g14387 ( n15964 , n19983 , n11577 );
    xnor g14388 ( n10674 , n12651 , n28612 );
    xnor g14389 ( n27718 , n2853 , n3846 );
    not g14390 ( n7670 , n8947 );
    or g14391 ( n7309 , n21725 , n6598 );
    nor g14392 ( n25886 , n14430 , n31513 );
    xnor g14393 ( n14602 , n4929 , n2483 );
    nor g14394 ( n1985 , n9336 , n6811 );
    or g14395 ( n5063 , n15989 , n20321 );
    or g14396 ( n8138 , n31133 , n24011 );
    not g14397 ( n1379 , n6254 );
    xor g14398 ( n30997 , n19427 , n20622 );
    xnor g14399 ( n9959 , n25715 , n28993 );
    not g14400 ( n22595 , n31889 );
    or g14401 ( n3018 , n27929 , n18525 );
    or g14402 ( n7831 , n5611 , n29178 );
    not g14403 ( n2568 , n754 );
    not g14404 ( n17391 , n20436 );
    not g14405 ( n18575 , n21107 );
    not g14406 ( n15335 , n17475 );
    or g14407 ( n23509 , n7404 , n12068 );
    and g14408 ( n19310 , n16687 , n5758 );
    or g14409 ( n22137 , n26052 , n13242 );
    xnor g14410 ( n10236 , n26550 , n14548 );
    or g14411 ( n7666 , n6456 , n27947 );
    or g14412 ( n27436 , n22808 , n31434 );
    nor g14413 ( n14493 , n1670 , n11392 );
    xnor g14414 ( n1810 , n10346 , n12312 );
    buf g14415 ( n30812 , n14854 );
    nor g14416 ( n19694 , n3036 , n31204 );
    xnor g14417 ( n16879 , n30580 , n14064 );
    not g14418 ( n7217 , n29148 );
    and g14419 ( n15323 , n24584 , n18004 );
    xnor g14420 ( n8754 , n27354 , n9619 );
    xnor g14421 ( n16329 , n25108 , n23796 );
    nor g14422 ( n17003 , n7855 , n26559 );
    not g14423 ( n21846 , n31785 );
    or g14424 ( n11567 , n24853 , n26945 );
    xor g14425 ( n20505 , n17060 , n3348 );
    and g14426 ( n21662 , n6790 , n20127 );
    or g14427 ( n26704 , n24218 , n3348 );
    or g14428 ( n14254 , n1635 , n9461 );
    and g14429 ( n761 , n668 , n25097 );
    and g14430 ( n30368 , n21188 , n23876 );
    not g14431 ( n12043 , n28281 );
    and g14432 ( n4355 , n30639 , n7377 );
    not g14433 ( n12341 , n12607 );
    not g14434 ( n29857 , n11804 );
    and g14435 ( n26887 , n17347 , n24066 );
    or g14436 ( n22477 , n24408 , n15054 );
    nor g14437 ( n8879 , n9163 , n12596 );
    buf g14438 ( n11313 , n22454 );
    or g14439 ( n30847 , n29604 , n18984 );
    xnor g14440 ( n8706 , n25964 , n31427 );
    xnor g14441 ( n6430 , n18456 , n18675 );
    and g14442 ( n8818 , n24447 , n2899 );
    xnor g14443 ( n2632 , n10768 , n27829 );
    or g14444 ( n9581 , n14400 , n3618 );
    not g14445 ( n1105 , n10853 );
    not g14446 ( n5979 , n16019 );
    and g14447 ( n12463 , n5658 , n17043 );
    xnor g14448 ( n6309 , n1315 , n26191 );
    or g14449 ( n1174 , n7368 , n22276 );
    xnor g14450 ( n16376 , n17771 , n4662 );
    xnor g14451 ( n15947 , n8659 , n27973 );
    or g14452 ( n27977 , n4582 , n10634 );
    not g14453 ( n24568 , n2548 );
    not g14454 ( n10203 , n25424 );
    not g14455 ( n5456 , n1635 );
    not g14456 ( n9894 , n21289 );
    not g14457 ( n22111 , n17563 );
    xnor g14458 ( n28389 , n16299 , n20198 );
    not g14459 ( n22401 , n11234 );
    nor g14460 ( n19454 , n4468 , n31691 );
    not g14461 ( n2511 , n11658 );
    xnor g14462 ( n7926 , n20226 , n793 );
    and g14463 ( n12719 , n20076 , n2930 );
    nor g14464 ( n17484 , n23634 , n13627 );
    not g14465 ( n24407 , n9822 );
    and g14466 ( n24140 , n18593 , n13019 );
    and g14467 ( n20449 , n27701 , n30471 );
    xor g14468 ( n20853 , n7661 , n25678 );
    not g14469 ( n24138 , n1432 );
    xnor g14470 ( n30412 , n30752 , n29667 );
    or g14471 ( n29799 , n421 , n21278 );
    xnor g14472 ( n1342 , n3073 , n12215 );
    and g14473 ( n17031 , n8343 , n24162 );
    or g14474 ( n4945 , n25143 , n25283 );
    xnor g14475 ( n17478 , n7618 , n5656 );
    not g14476 ( n6464 , n12897 );
    or g14477 ( n28421 , n9866 , n14461 );
    not g14478 ( n31196 , n13454 );
    or g14479 ( n8060 , n30804 , n18703 );
    and g14480 ( n29357 , n12099 , n10643 );
    xnor g14481 ( n31842 , n8929 , n14145 );
    and g14482 ( n27795 , n29429 , n10547 );
    xnor g14483 ( n6253 , n7061 , n1495 );
    xnor g14484 ( n14069 , n10827 , n8834 );
    xnor g14485 ( n25947 , n11603 , n26062 );
    nor g14486 ( n29216 , n8893 , n27345 );
    nor g14487 ( n31703 , n20750 , n19726 );
    and g14488 ( n13322 , n1155 , n28228 );
    not g14489 ( n31230 , n31821 );
    xnor g14490 ( n32032 , n1460 , n23514 );
    xnor g14491 ( n8088 , n2473 , n18612 );
    or g14492 ( n4470 , n18667 , n17904 );
    not g14493 ( n19683 , n15211 );
    not g14494 ( n5489 , n14123 );
    and g14495 ( n13156 , n28846 , n27843 );
    xnor g14496 ( n18100 , n26363 , n4988 );
    xnor g14497 ( n4533 , n30459 , n14400 );
    not g14498 ( n4260 , n17912 );
    not g14499 ( n11594 , n2190 );
    or g14500 ( n31251 , n16721 , n23815 );
    xnor g14501 ( n20722 , n11352 , n4503 );
    nor g14502 ( n15632 , n4339 , n24445 );
    not g14503 ( n3689 , n4796 );
    nor g14504 ( n2763 , n22922 , n3933 );
    and g14505 ( n26194 , n14938 , n8943 );
    or g14506 ( n18777 , n24948 , n19117 );
    nor g14507 ( n25236 , n26002 , n1095 );
    xnor g14508 ( n28270 , n1586 , n27562 );
    not g14509 ( n18893 , n25146 );
    xnor g14510 ( n6660 , n13714 , n6223 );
    not g14511 ( n7748 , n31486 );
    not g14512 ( n27854 , n14387 );
    or g14513 ( n9662 , n19269 , n27751 );
    or g14514 ( n18864 , n22206 , n7865 );
    or g14515 ( n18591 , n7598 , n27635 );
    not g14516 ( n18975 , n30497 );
    or g14517 ( n4395 , n28341 , n4246 );
    and g14518 ( n23315 , n26543 , n17964 );
    xnor g14519 ( n30477 , n11361 , n6306 );
    not g14520 ( n3845 , n30982 );
    xor g14521 ( n15534 , n11901 , n30510 );
    xnor g14522 ( n10852 , n28734 , n28562 );
    and g14523 ( n9210 , n7509 , n18814 );
    and g14524 ( n24555 , n12981 , n20814 );
    xnor g14525 ( n10251 , n13954 , n28046 );
    and g14526 ( n24001 , n21203 , n11356 );
    or g14527 ( n7236 , n2856 , n969 );
    not g14528 ( n6194 , n13332 );
    and g14529 ( n17541 , n4198 , n24531 );
    xnor g14530 ( n7668 , n17719 , n20763 );
    nor g14531 ( n81 , n28911 , n14770 );
    not g14532 ( n4624 , n6533 );
    xnor g14533 ( n2552 , n19286 , n5449 );
    or g14534 ( n20496 , n10924 , n22639 );
    or g14535 ( n18594 , n25094 , n30362 );
    not g14536 ( n11381 , n1127 );
    or g14537 ( n7211 , n1091 , n23850 );
    xnor g14538 ( n7708 , n25598 , n6099 );
    xnor g14539 ( n2836 , n30671 , n31482 );
    and g14540 ( n30804 , n7857 , n19300 );
    not g14541 ( n22264 , n24676 );
    not g14542 ( n8198 , n4351 );
    xnor g14543 ( n3241 , n19758 , n12363 );
    not g14544 ( n3763 , n947 );
    and g14545 ( n14717 , n14722 , n16049 );
    not g14546 ( n6162 , n2071 );
    not g14547 ( n14332 , n13734 );
    not g14548 ( n13467 , n2212 );
    not g14549 ( n15819 , n15987 );
    or g14550 ( n27479 , n15119 , n19686 );
    xnor g14551 ( n8787 , n29782 , n24386 );
    xnor g14552 ( n20846 , n11004 , n24107 );
    and g14553 ( n18115 , n12472 , n5996 );
    and g14554 ( n5520 , n20530 , n16078 );
    and g14555 ( n31247 , n20912 , n613 );
    or g14556 ( n17306 , n2273 , n2983 );
    xnor g14557 ( n6354 , n12537 , n6138 );
    not g14558 ( n4735 , n9865 );
    nor g14559 ( n4941 , n22217 , n24979 );
    or g14560 ( n1124 , n11281 , n6937 );
    xnor g14561 ( n31453 , n13463 , n24949 );
    and g14562 ( n29754 , n25873 , n27516 );
    xnor g14563 ( n17316 , n10778 , n14398 );
    and g14564 ( n31121 , n14939 , n20978 );
    not g14565 ( n22692 , n8443 );
    or g14566 ( n26199 , n2963 , n25069 );
    not g14567 ( n2834 , n18404 );
    xnor g14568 ( n15124 , n15235 , n13936 );
    and g14569 ( n19303 , n11093 , n11723 );
    not g14570 ( n4946 , n20041 );
    or g14571 ( n24779 , n11535 , n15587 );
    or g14572 ( n3952 , n930 , n13441 );
    not g14573 ( n13585 , n17180 );
    xnor g14574 ( n6169 , n14795 , n18203 );
    xor g14575 ( n11860 , n31892 , n22296 );
    not g14576 ( n2317 , n22632 );
    not g14577 ( n21164 , n12866 );
    xor g14578 ( n26324 , n22041 , n9183 );
    xnor g14579 ( n18487 , n16576 , n23706 );
    xnor g14580 ( n2740 , n25363 , n12715 );
    and g14581 ( n28126 , n31571 , n6916 );
    xnor g14582 ( n21614 , n21273 , n15842 );
    xnor g14583 ( n26549 , n26013 , n26462 );
    xor g14584 ( n7109 , n28412 , n25672 );
    not g14585 ( n24596 , n5518 );
    not g14586 ( n31667 , n23045 );
    nor g14587 ( n28926 , n22415 , n11552 );
    and g14588 ( n29340 , n28307 , n5945 );
    not g14589 ( n31526 , n20955 );
    buf g14590 ( n4632 , n9418 );
    or g14591 ( n7056 , n21383 , n27538 );
    not g14592 ( n21534 , n12756 );
    and g14593 ( n4206 , n10780 , n2811 );
    nor g14594 ( n9969 , n24607 , n16054 );
    or g14595 ( n9398 , n2326 , n12629 );
    nor g14596 ( n1359 , n793 , n5386 );
    and g14597 ( n29614 , n25588 , n10895 );
    xnor g14598 ( n10506 , n31222 , n23064 );
    not g14599 ( n2541 , n22450 );
    not g14600 ( n29584 , n10367 );
    xnor g14601 ( n9141 , n6299 , n27988 );
    xnor g14602 ( n7138 , n26697 , n16204 );
    or g14603 ( n18673 , n15082 , n14506 );
    xnor g14604 ( n12472 , n8276 , n24714 );
    not g14605 ( n28156 , n5982 );
    and g14606 ( n279 , n1619 , n25521 );
    or g14607 ( n28730 , n9765 , n20010 );
    or g14608 ( n7544 , n31850 , n26471 );
    not g14609 ( n23928 , n7439 );
    nor g14610 ( n19076 , n2078 , n27272 );
    xnor g14611 ( n23752 , n14898 , n13059 );
    or g14612 ( n20500 , n12585 , n23854 );
    not g14613 ( n16248 , n6419 );
    and g14614 ( n2285 , n26990 , n27494 );
    not g14615 ( n4623 , n30256 );
    not g14616 ( n9541 , n30790 );
    xnor g14617 ( n15804 , n30527 , n4472 );
    xnor g14618 ( n4177 , n2767 , n26581 );
    not g14619 ( n4087 , n7717 );
    and g14620 ( n19890 , n12378 , n2453 );
    xnor g14621 ( n19654 , n9222 , n2986 );
    not g14622 ( n3483 , n1815 );
    not g14623 ( n6325 , n7157 );
    nor g14624 ( n27573 , n19945 , n6159 );
    or g14625 ( n18268 , n20646 , n25352 );
    or g14626 ( n13856 , n27674 , n11656 );
    not g14627 ( n3077 , n19924 );
    not g14628 ( n4252 , n19328 );
    not g14629 ( n2801 , n24540 );
    not g14630 ( n20823 , n28931 );
    nor g14631 ( n19507 , n3706 , n3427 );
    or g14632 ( n31135 , n19665 , n28652 );
    not g14633 ( n15676 , n22854 );
    xnor g14634 ( n2092 , n8603 , n13177 );
    not g14635 ( n17435 , n27144 );
    not g14636 ( n6251 , n13325 );
    or g14637 ( n23916 , n31808 , n13650 );
    and g14638 ( n7273 , n9268 , n21046 );
    and g14639 ( n15921 , n18228 , n7040 );
    not g14640 ( n27842 , n18995 );
    xnor g14641 ( n12338 , n19267 , n12347 );
    and g14642 ( n18337 , n1038 , n24701 );
    not g14643 ( n19326 , n26758 );
    not g14644 ( n15734 , n5251 );
    xor g14645 ( n1425 , n31472 , n12518 );
    and g14646 ( n12316 , n30003 , n19700 );
    nor g14647 ( n22602 , n16540 , n15934 );
    xnor g14648 ( n25024 , n5171 , n31088 );
    not g14649 ( n652 , n30006 );
    not g14650 ( n22897 , n11039 );
    not g14651 ( n15192 , n24164 );
    xor g14652 ( n17763 , n4700 , n1095 );
    or g14653 ( n10221 , n27627 , n7481 );
    not g14654 ( n18198 , n27637 );
    or g14655 ( n2152 , n2872 , n18783 );
    xnor g14656 ( n8915 , n24197 , n30214 );
    xor g14657 ( n28046 , n12964 , n20870 );
    or g14658 ( n127 , n14393 , n3838 );
    and g14659 ( n8175 , n23219 , n7994 );
    and g14660 ( n4528 , n542 , n7884 );
    xnor g14661 ( n5330 , n8698 , n17782 );
    or g14662 ( n12724 , n21720 , n24981 );
    not g14663 ( n26436 , n16991 );
    xnor g14664 ( n10263 , n29482 , n1760 );
    nor g14665 ( n26155 , n12612 , n21175 );
    xnor g14666 ( n22798 , n3997 , n12263 );
    xnor g14667 ( n17427 , n3920 , n13663 );
    or g14668 ( n16541 , n14805 , n27264 );
    and g14669 ( n30919 , n14485 , n1384 );
    not g14670 ( n30389 , n980 );
    or g14671 ( n15263 , n8869 , n30820 );
    xnor g14672 ( n21033 , n3790 , n24182 );
    or g14673 ( n6198 , n3654 , n28859 );
    or g14674 ( n24299 , n10139 , n3799 );
    xnor g14675 ( n20874 , n528 , n28305 );
    or g14676 ( n12421 , n4463 , n4478 );
    and g14677 ( n12828 , n6279 , n27608 );
    not g14678 ( n17248 , n17255 );
    and g14679 ( n27173 , n19387 , n24098 );
    not g14680 ( n23358 , n9434 );
    not g14681 ( n28904 , n14136 );
    or g14682 ( n14682 , n19168 , n24062 );
    xnor g14683 ( n10686 , n9189 , n1020 );
    not g14684 ( n19687 , n9509 );
    xnor g14685 ( n3254 , n20698 , n11643 );
    or g14686 ( n11455 , n20623 , n11033 );
    xnor g14687 ( n24626 , n15091 , n21716 );
    not g14688 ( n23819 , n29407 );
    xnor g14689 ( n25768 , n11824 , n13357 );
    and g14690 ( n26733 , n7894 , n20366 );
    xnor g14691 ( n8513 , n13396 , n6310 );
    or g14692 ( n17485 , n13859 , n15214 );
    not g14693 ( n30481 , n21977 );
    and g14694 ( n7328 , n30070 , n7773 );
    xnor g14695 ( n17902 , n29749 , n23694 );
    not g14696 ( n6676 , n4298 );
    xnor g14697 ( n28830 , n23456 , n23681 );
    not g14698 ( n30866 , n21442 );
    xnor g14699 ( n25065 , n31773 , n9653 );
    not g14700 ( n29108 , n19679 );
    not g14701 ( n7349 , n16448 );
    or g14702 ( n9344 , n18871 , n12273 );
    not g14703 ( n23585 , n4096 );
    xnor g14704 ( n27252 , n31936 , n14599 );
    xnor g14705 ( n15484 , n22438 , n13612 );
    or g14706 ( n31903 , n25773 , n19585 );
    or g14707 ( n27111 , n14566 , n17313 );
    xnor g14708 ( n22954 , n29231 , n30063 );
    xnor g14709 ( n29086 , n8815 , n15210 );
    xnor g14710 ( n12729 , n24935 , n20067 );
    xnor g14711 ( n25448 , n31041 , n7080 );
    xnor g14712 ( n15849 , n1907 , n9439 );
    or g14713 ( n30589 , n18045 , n21107 );
    xnor g14714 ( n1213 , n19354 , n17771 );
    not g14715 ( n6904 , n11743 );
    or g14716 ( n25609 , n30947 , n29449 );
    nor g14717 ( n26540 , n15977 , n12188 );
    xnor g14718 ( n19477 , n30436 , n30378 );
    xnor g14719 ( n21880 , n19641 , n15191 );
    and g14720 ( n20465 , n12890 , n3000 );
    not g14721 ( n12760 , n22905 );
    not g14722 ( n14539 , n24271 );
    nor g14723 ( n22427 , n11643 , n31070 );
    nor g14724 ( n27247 , n25842 , n19157 );
    not g14725 ( n203 , n1524 );
    nor g14726 ( n1153 , n20486 , n11523 );
    xnor g14727 ( n11346 , n14518 , n320 );
    or g14728 ( n3922 , n29632 , n14249 );
    or g14729 ( n13080 , n7473 , n5677 );
    or g14730 ( n19307 , n11019 , n18430 );
    xnor g14731 ( n17312 , n4939 , n23115 );
    or g14732 ( n1227 , n8986 , n1204 );
    and g14733 ( n16555 , n8160 , n18641 );
    or g14734 ( n26450 , n4352 , n17618 );
    or g14735 ( n24805 , n29090 , n813 );
    xor g14736 ( n14826 , n12505 , n19889 );
    and g14737 ( n5363 , n28377 , n14581 );
    not g14738 ( n259 , n5012 );
    not g14739 ( n13441 , n19600 );
    xnor g14740 ( n10868 , n860 , n5944 );
    not g14741 ( n12285 , n554 );
    xnor g14742 ( n11488 , n8079 , n5457 );
    and g14743 ( n24627 , n10757 , n11032 );
    xnor g14744 ( n25396 , n20520 , n9746 );
    xnor g14745 ( n21359 , n16429 , n23748 );
    and g14746 ( n11042 , n3024 , n22128 );
    or g14747 ( n23214 , n17551 , n3662 );
    and g14748 ( n26818 , n3899 , n17105 );
    not g14749 ( n10738 , n5930 );
    xnor g14750 ( n26752 , n21064 , n19632 );
    xnor g14751 ( n2559 , n22132 , n8797 );
    xnor g14752 ( n6371 , n15426 , n31933 );
    nor g14753 ( n18838 , n24132 , n12652 );
    nor g14754 ( n2716 , n27453 , n31896 );
    or g14755 ( n23860 , n8313 , n24135 );
    nor g14756 ( n7175 , n19575 , n18671 );
    or g14757 ( n12303 , n16135 , n13032 );
    not g14758 ( n14447 , n1027 );
    or g14759 ( n12981 , n23522 , n5462 );
    and g14760 ( n25578 , n20974 , n23352 );
    not g14761 ( n15557 , n10034 );
    not g14762 ( n11309 , n21701 );
    and g14763 ( n102 , n15451 , n29853 );
    or g14764 ( n15284 , n11581 , n17376 );
    and g14765 ( n6982 , n6545 , n24312 );
    or g14766 ( n3966 , n14452 , n6284 );
    xnor g14767 ( n24974 , n11104 , n25219 );
    not g14768 ( n10179 , n20476 );
    not g14769 ( n2539 , n24794 );
    and g14770 ( n20219 , n9641 , n12417 );
    xnor g14771 ( n24238 , n31059 , n3621 );
    nor g14772 ( n13736 , n22073 , n21182 );
    and g14773 ( n20809 , n22989 , n20635 );
    and g14774 ( n19007 , n443 , n23169 );
    and g14775 ( n14304 , n2367 , n9360 );
    or g14776 ( n8113 , n6211 , n18139 );
    xnor g14777 ( n25774 , n14740 , n25446 );
    or g14778 ( n20362 , n3570 , n25935 );
    xnor g14779 ( n30275 , n15090 , n29818 );
    not g14780 ( n9446 , n10777 );
    not g14781 ( n9473 , n13571 );
    xnor g14782 ( n14623 , n8708 , n26226 );
    not g14783 ( n27438 , n20080 );
    not g14784 ( n7438 , n10802 );
    not g14785 ( n8956 , n12900 );
    or g14786 ( n26739 , n3591 , n15663 );
    nor g14787 ( n22536 , n13415 , n547 );
    xnor g14788 ( n5690 , n31061 , n22037 );
    not g14789 ( n24788 , n19462 );
    xnor g14790 ( n7698 , n23173 , n27672 );
    not g14791 ( n28133 , n10784 );
    xnor g14792 ( n23198 , n20680 , n2862 );
    xnor g14793 ( n1255 , n18709 , n28799 );
    xnor g14794 ( n18986 , n21618 , n24633 );
    xnor g14795 ( n20337 , n4490 , n26920 );
    and g14796 ( n28866 , n25340 , n8096 );
    nor g14797 ( n338 , n16908 , n9983 );
    or g14798 ( n12314 , n24351 , n31101 );
    and g14799 ( n22943 , n19437 , n16161 );
    xnor g14800 ( n10680 , n17893 , n22244 );
    and g14801 ( n4563 , n1876 , n20626 );
    xnor g14802 ( n29363 , n24045 , n21680 );
    not g14803 ( n17016 , n20051 );
    not g14804 ( n26208 , n6076 );
    not g14805 ( n10818 , n30209 );
    or g14806 ( n26154 , n2453 , n12378 );
    xnor g14807 ( n23317 , n1568 , n22178 );
    xnor g14808 ( n22679 , n9145 , n7787 );
    not g14809 ( n30596 , n17793 );
    not g14810 ( n23380 , n25860 );
    or g14811 ( n29704 , n11058 , n28839 );
    not g14812 ( n8774 , n22094 );
    xnor g14813 ( n9277 , n25954 , n2748 );
    not g14814 ( n11693 , n2095 );
    and g14815 ( n26810 , n25845 , n23570 );
    not g14816 ( n4151 , n29673 );
    or g14817 ( n22853 , n19103 , n537 );
    or g14818 ( n8864 , n27034 , n8436 );
    xnor g14819 ( n29718 , n19231 , n4358 );
    nor g14820 ( n6987 , n14093 , n26768 );
    or g14821 ( n7038 , n6196 , n18504 );
    xnor g14822 ( n28032 , n6777 , n3376 );
    xnor g14823 ( n31299 , n25893 , n25546 );
    not g14824 ( n9461 , n3432 );
    and g14825 ( n10546 , n18026 , n1035 );
    not g14826 ( n3744 , n18199 );
    not g14827 ( n15948 , n11360 );
    xnor g14828 ( n1781 , n2243 , n6482 );
    and g14829 ( n15925 , n14334 , n15911 );
    not g14830 ( n11660 , n54 );
    nor g14831 ( n14871 , n22248 , n12990 );
    nor g14832 ( n18733 , n23960 , n23647 );
    xnor g14833 ( n3916 , n16459 , n18203 );
    xnor g14834 ( n21921 , n20502 , n16529 );
    or g14835 ( n24842 , n7345 , n25212 );
    xnor g14836 ( n24820 , n19716 , n20510 );
    or g14837 ( n3217 , n6151 , n18961 );
    xnor g14838 ( n15499 , n19877 , n17236 );
    not g14839 ( n9809 , n30069 );
    xnor g14840 ( n13964 , n24592 , n19574 );
    not g14841 ( n920 , n9087 );
    xnor g14842 ( n2069 , n18074 , n9529 );
    or g14843 ( n30810 , n22165 , n1187 );
    and g14844 ( n11923 , n16067 , n29385 );
    not g14845 ( n7431 , n25136 );
    not g14846 ( n12859 , n26162 );
    xnor g14847 ( n24561 , n24418 , n20825 );
    and g14848 ( n22755 , n25409 , n11680 );
    and g14849 ( n21111 , n23479 , n20119 );
    or g14850 ( n20541 , n1846 , n8863 );
    xnor g14851 ( n583 , n24660 , n3059 );
    nor g14852 ( n7533 , n7655 , n3787 );
    or g14853 ( n27144 , n1616 , n20754 );
    xnor g14854 ( n28098 , n30146 , n31829 );
    nor g14855 ( n5607 , n7539 , n6162 );
    not g14856 ( n735 , n22844 );
    or g14857 ( n16226 , n10997 , n21769 );
    or g14858 ( n13272 , n489 , n8349 );
    not g14859 ( n26666 , n12321 );
    xnor g14860 ( n20653 , n22441 , n8005 );
    not g14861 ( n19069 , n6435 );
    not g14862 ( n7930 , n28325 );
    not g14863 ( n5006 , n28378 );
    or g14864 ( n29624 , n22240 , n3183 );
    and g14865 ( n28442 , n16886 , n19455 );
    xnor g14866 ( n13895 , n3116 , n7969 );
    not g14867 ( n19734 , n8623 );
    xnor g14868 ( n707 , n25563 , n8713 );
    xnor g14869 ( n21125 , n27297 , n7107 );
    not g14870 ( n18410 , n9301 );
    xnor g14871 ( n19038 , n17068 , n6349 );
    or g14872 ( n9603 , n9520 , n20334 );
    nor g14873 ( n18342 , n13137 , n27805 );
    and g14874 ( n22860 , n1583 , n11978 );
    not g14875 ( n5543 , n25978 );
    nor g14876 ( n31589 , n29601 , n4682 );
    or g14877 ( n18445 , n5857 , n19724 );
    not g14878 ( n9710 , n15181 );
    not g14879 ( n14517 , n8742 );
    not g14880 ( n16535 , n28808 );
    or g14881 ( n4597 , n11119 , n28487 );
    or g14882 ( n14007 , n16572 , n17512 );
    or g14883 ( n27683 , n19694 , n25377 );
    xnor g14884 ( n7878 , n17810 , n26246 );
    not g14885 ( n18502 , n11098 );
    and g14886 ( n17926 , n5676 , n15222 );
    nor g14887 ( n19849 , n3725 , n21709 );
    nor g14888 ( n8464 , n13317 , n24241 );
    xnor g14889 ( n3843 , n9586 , n7740 );
    or g14890 ( n23977 , n8683 , n31552 );
    and g14891 ( n136 , n7856 , n2816 );
    or g14892 ( n23821 , n2037 , n13926 );
    nor g14893 ( n9559 , n22922 , n12159 );
    or g14894 ( n7468 , n21104 , n25791 );
    and g14895 ( n28107 , n20872 , n8390 );
    or g14896 ( n491 , n16439 , n28639 );
    nor g14897 ( n31107 , n19790 , n27058 );
    not g14898 ( n5729 , n17295 );
    not g14899 ( n29170 , n18184 );
    not g14900 ( n25981 , n11847 );
    or g14901 ( n20136 , n12050 , n25918 );
    nor g14902 ( n26504 , n17983 , n18143 );
    or g14903 ( n1877 , n2414 , n3457 );
    xnor g14904 ( n8001 , n12406 , n31224 );
    xnor g14905 ( n7795 , n26899 , n5734 );
    not g14906 ( n5996 , n15417 );
    and g14907 ( n2544 , n31890 , n3837 );
    xnor g14908 ( n1406 , n25025 , n10177 );
    and g14909 ( n2321 , n7869 , n15902 );
    xor g14910 ( n26418 , n1803 , n13298 );
    or g14911 ( n6239 , n25284 , n11305 );
    xnor g14912 ( n3346 , n291 , n30321 );
    xnor g14913 ( n30823 , n5360 , n13640 );
    not g14914 ( n25395 , n11491 );
    xnor g14915 ( n7110 , n26340 , n22751 );
    xor g14916 ( n121 , n16857 , n14246 );
    xnor g14917 ( n21312 , n11569 , n31124 );
    and g14918 ( n9462 , n17553 , n27592 );
    xnor g14919 ( n15040 , n12434 , n4421 );
    or g14920 ( n10809 , n5876 , n19790 );
    xnor g14921 ( n22411 , n7419 , n4020 );
    or g14922 ( n14501 , n30574 , n4949 );
    and g14923 ( n4441 , n13511 , n10798 );
    xnor g14924 ( n16765 , n9604 , n16998 );
    and g14925 ( n19818 , n6742 , n11236 );
    nor g14926 ( n5900 , n24230 , n7524 );
    and g14927 ( n20731 , n13537 , n27912 );
    or g14928 ( n8951 , n7613 , n23220 );
    xnor g14929 ( n26368 , n2926 , n13016 );
    not g14930 ( n10662 , n29845 );
    xnor g14931 ( n1733 , n18311 , n4149 );
    not g14932 ( n14039 , n8260 );
    nor g14933 ( n1597 , n10634 , n23050 );
    not g14934 ( n20803 , n30786 );
    or g14935 ( n25697 , n16435 , n9677 );
    or g14936 ( n9394 , n27286 , n19111 );
    nor g14937 ( n3357 , n9604 , n16998 );
    or g14938 ( n3495 , n17446 , n11818 );
    not g14939 ( n21616 , n8558 );
    nor g14940 ( n5431 , n6721 , n26505 );
    not g14941 ( n11205 , n12057 );
    not g14942 ( n15862 , n26690 );
    or g14943 ( n2891 , n26598 , n17506 );
    not g14944 ( n483 , n28183 );
    not g14945 ( n8726 , n18700 );
    not g14946 ( n28894 , n27868 );
    or g14947 ( n8494 , n26726 , n2082 );
    and g14948 ( n30527 , n7364 , n13740 );
    not g14949 ( n4619 , n21185 );
    or g14950 ( n2962 , n8988 , n20186 );
    and g14951 ( n10607 , n18844 , n923 );
    xnor g14952 ( n24134 , n2759 , n5708 );
    not g14953 ( n21736 , n16835 );
    and g14954 ( n6094 , n16141 , n10704 );
    or g14955 ( n21294 , n11905 , n14629 );
    not g14956 ( n30695 , n17195 );
    and g14957 ( n19760 , n2594 , n27451 );
    xnor g14958 ( n12554 , n3512 , n30717 );
    not g14959 ( n6500 , n29192 );
    not g14960 ( n901 , n21342 );
    xnor g14961 ( n22241 , n28382 , n1043 );
    xnor g14962 ( n10866 , n5092 , n20075 );
    not g14963 ( n22450 , n18821 );
    xnor g14964 ( n5515 , n11736 , n4213 );
    not g14965 ( n27635 , n327 );
    xnor g14966 ( n31464 , n29335 , n27885 );
    not g14967 ( n4686 , n16053 );
    and g14968 ( n2369 , n26528 , n24533 );
    xnor g14969 ( n2061 , n11309 , n15056 );
    or g14970 ( n1992 , n21564 , n8906 );
    nor g14971 ( n10369 , n19632 , n4004 );
    xnor g14972 ( n11940 , n19830 , n12821 );
    xnor g14973 ( n13179 , n14138 , n18683 );
    and g14974 ( n24923 , n23988 , n20963 );
    xnor g14975 ( n2535 , n29430 , n10158 );
    and g14976 ( n24806 , n19116 , n24772 );
    and g14977 ( n23128 , n30332 , n2812 );
    not g14978 ( n31930 , n26758 );
    not g14979 ( n21105 , n17019 );
    nor g14980 ( n18785 , n25391 , n20543 );
    xor g14981 ( n5656 , n3747 , n5638 );
    xnor g14982 ( n28090 , n25268 , n15226 );
    or g14983 ( n9320 , n25874 , n10793 );
    or g14984 ( n11762 , n3588 , n21292 );
    not g14985 ( n4862 , n19783 );
    xnor g14986 ( n20213 , n13119 , n3370 );
    nor g14987 ( n398 , n15258 , n12385 );
    or g14988 ( n1922 , n24840 , n13651 );
    or g14989 ( n9970 , n27805 , n15730 );
    not g14990 ( n15997 , n124 );
    and g14991 ( n25918 , n2158 , n29396 );
    not g14992 ( n12802 , n21585 );
    or g14993 ( n8500 , n23978 , n16859 );
    not g14994 ( n28150 , n29741 );
    nor g14995 ( n22126 , n6432 , n20280 );
    xnor g14996 ( n5593 , n18437 , n23740 );
    nor g14997 ( n16626 , n2453 , n20856 );
    and g14998 ( n3053 , n23930 , n21635 );
    not g14999 ( n4040 , n17998 );
    or g15000 ( n25961 , n9005 , n25946 );
    xor g15001 ( n6848 , n16274 , n27373 );
    not g15002 ( n27186 , n9098 );
    not g15003 ( n25610 , n4222 );
    and g15004 ( n21674 , n21715 , n648 );
    xnor g15005 ( n23516 , n23274 , n31620 );
    or g15006 ( n7463 , n6368 , n27599 );
    xnor g15007 ( n19433 , n23880 , n22389 );
    nor g15008 ( n21604 , n6509 , n30896 );
    or g15009 ( n17434 , n7156 , n5397 );
    and g15010 ( n5892 , n28857 , n6603 );
    or g15011 ( n29752 , n8306 , n28152 );
    or g15012 ( n24708 , n31056 , n14097 );
    or g15013 ( n23482 , n24404 , n3986 );
    and g15014 ( n7222 , n6908 , n26597 );
    or g15015 ( n28343 , n21621 , n17018 );
    and g15016 ( n16317 , n214 , n15737 );
    not g15017 ( n23176 , n3131 );
    nor g15018 ( n19166 , n22259 , n16133 );
    and g15019 ( n3239 , n28929 , n14693 );
    and g15020 ( n14020 , n28714 , n3809 );
    or g15021 ( n23498 , n26116 , n582 );
    or g15022 ( n1074 , n3081 , n4983 );
    or g15023 ( n6001 , n4057 , n21932 );
    not g15024 ( n29016 , n15733 );
    not g15025 ( n17521 , n30806 );
    or g15026 ( n30070 , n20356 , n14799 );
    xnor g15027 ( n17329 , n29642 , n5521 );
    and g15028 ( n27219 , n14394 , n25466 );
    xnor g15029 ( n21139 , n12598 , n28441 );
    and g15030 ( n30047 , n19155 , n13140 );
    and g15031 ( n5759 , n16148 , n22881 );
    and g15032 ( n25831 , n10033 , n4217 );
    nor g15033 ( n1247 , n3360 , n26644 );
    or g15034 ( n10632 , n21508 , n8870 );
    and g15035 ( n5440 , n28314 , n12035 );
    or g15036 ( n1594 , n28680 , n20992 );
    not g15037 ( n11706 , n18199 );
    and g15038 ( n15668 , n16232 , n4011 );
    xnor g15039 ( n15886 , n14275 , n8118 );
    not g15040 ( n3315 , n22174 );
    nor g15041 ( n8521 , n31676 , n26373 );
    buf g15042 ( n6071 , n22620 );
    not g15043 ( n3797 , n977 );
    not g15044 ( n19865 , n13225 );
    xnor g15045 ( n11679 , n16056 , n2487 );
    or g15046 ( n26222 , n25472 , n18789 );
    nor g15047 ( n22487 , n3108 , n29552 );
    xnor g15048 ( n29014 , n16799 , n26114 );
    xnor g15049 ( n28216 , n28305 , n350 );
    or g15050 ( n30808 , n1464 , n6876 );
    nor g15051 ( n31184 , n25971 , n4474 );
    nor g15052 ( n9598 , n1692 , n21023 );
    not g15053 ( n15276 , n14800 );
    not g15054 ( n30522 , n1477 );
    xnor g15055 ( n31427 , n15525 , n17775 );
    xnor g15056 ( n12063 , n28470 , n31889 );
    or g15057 ( n13605 , n27930 , n19042 );
    or g15058 ( n25052 , n29574 , n13086 );
    or g15059 ( n14781 , n27011 , n29 );
    or g15060 ( n9993 , n18455 , n20172 );
    not g15061 ( n7604 , n30490 );
    or g15062 ( n1911 , n7836 , n23973 );
    not g15063 ( n18775 , n25387 );
    xnor g15064 ( n27153 , n28693 , n7513 );
    nor g15065 ( n295 , n12221 , n13836 );
    xnor g15066 ( n26778 , n29894 , n15463 );
    not g15067 ( n14238 , n13285 );
    or g15068 ( n2458 , n12550 , n5895 );
    xnor g15069 ( n24050 , n26052 , n2001 );
    xnor g15070 ( n14073 , n23526 , n10319 );
    nor g15071 ( n5952 , n22549 , n608 );
    xnor g15072 ( n11948 , n12399 , n7473 );
    not g15073 ( n8450 , n27064 );
    or g15074 ( n18964 , n31819 , n5322 );
    not g15075 ( n19617 , n28837 );
    not g15076 ( n17506 , n11060 );
    and g15077 ( n16153 , n1517 , n24509 );
    xnor g15078 ( n11547 , n22893 , n31473 );
    xnor g15079 ( n27325 , n20313 , n3080 );
    and g15080 ( n18715 , n12198 , n19217 );
    not g15081 ( n25893 , n17112 );
    not g15082 ( n1471 , n18504 );
    not g15083 ( n18997 , n13698 );
    not g15084 ( n11159 , n26585 );
    xnor g15085 ( n1567 , n16695 , n11343 );
    xnor g15086 ( n19067 , n27604 , n7931 );
    xnor g15087 ( n25048 , n18655 , n26398 );
    xnor g15088 ( n23568 , n4466 , n22045 );
    xnor g15089 ( n27752 , n3275 , n6135 );
    or g15090 ( n14746 , n13604 , n30290 );
    not g15091 ( n28044 , n26091 );
    not g15092 ( n10068 , n7209 );
    and g15093 ( n28197 , n5370 , n4871 );
    xnor g15094 ( n11921 , n17256 , n4324 );
    and g15095 ( n31499 , n1218 , n2684 );
    xnor g15096 ( n2829 , n31216 , n14109 );
    or g15097 ( n21548 , n19745 , n30783 );
    and g15098 ( n26950 , n30852 , n18398 );
    not g15099 ( n4749 , n23246 );
    nor g15100 ( n6271 , n17851 , n2618 );
    or g15101 ( n19991 , n16147 , n25590 );
    or g15102 ( n10184 , n24660 , n3059 );
    nor g15103 ( n9876 , n12364 , n13840 );
    xnor g15104 ( n20695 , n11335 , n26248 );
    or g15105 ( n18708 , n25933 , n31495 );
    nor g15106 ( n6807 , n7787 , n28694 );
    or g15107 ( n28508 , n11593 , n10030 );
    xnor g15108 ( n1881 , n15459 , n23613 );
    or g15109 ( n2322 , n30963 , n3893 );
    xnor g15110 ( n17354 , n17502 , n28963 );
    xnor g15111 ( n5254 , n24383 , n17126 );
    xnor g15112 ( n18542 , n24788 , n23232 );
    and g15113 ( n22374 , n27190 , n20506 );
    not g15114 ( n19886 , n17482 );
    xnor g15115 ( n24193 , n24585 , n8404 );
    xnor g15116 ( n15693 , n25283 , n29545 );
    and g15117 ( n26270 , n29219 , n4328 );
    xnor g15118 ( n15035 , n21601 , n24822 );
    not g15119 ( n11777 , n4663 );
    or g15120 ( n28771 , n26867 , n11484 );
    and g15121 ( n15646 , n12476 , n29652 );
    or g15122 ( n22265 , n24636 , n7181 );
    not g15123 ( n23549 , n15666 );
    not g15124 ( n24896 , n15122 );
    or g15125 ( n26871 , n2385 , n29515 );
    xnor g15126 ( n20019 , n16022 , n16788 );
    xnor g15127 ( n23800 , n6457 , n31267 );
    and g15128 ( n14250 , n6075 , n464 );
    or g15129 ( n2865 , n12637 , n26164 );
    not g15130 ( n3986 , n12964 );
    or g15131 ( n25151 , n2969 , n3055 );
    or g15132 ( n23020 , n23040 , n2939 );
    xnor g15133 ( n12938 , n6730 , n1565 );
    not g15134 ( n14657 , n11389 );
    not g15135 ( n20215 , n15710 );
    not g15136 ( n22136 , n5697 );
    or g15137 ( n3957 , n19190 , n2198 );
    xnor g15138 ( n17060 , n3943 , n30664 );
    and g15139 ( n10576 , n28194 , n31108 );
    and g15140 ( n8396 , n25321 , n27845 );
    and g15141 ( n31840 , n18926 , n31708 );
    not g15142 ( n11419 , n5521 );
    xnor g15143 ( n7187 , n14224 , n8094 );
    xnor g15144 ( n9369 , n2876 , n1381 );
    not g15145 ( n27330 , n16821 );
    not g15146 ( n28419 , n8031 );
    xnor g15147 ( n3084 , n9618 , n9062 );
    xnor g15148 ( n3179 , n15597 , n16551 );
    nor g15149 ( n15853 , n26941 , n3283 );
    xnor g15150 ( n25326 , n5364 , n11194 );
    not g15151 ( n27018 , n19879 );
    nor g15152 ( n13347 , n5361 , n17511 );
    xnor g15153 ( n17196 , n30983 , n7812 );
    nor g15154 ( n8546 , n25745 , n10853 );
    xnor g15155 ( n462 , n25765 , n26996 );
    not g15156 ( n19243 , n2566 );
    nor g15157 ( n4345 , n385 , n28028 );
    xnor g15158 ( n16180 , n13957 , n19300 );
    not g15159 ( n31131 , n14800 );
    or g15160 ( n15614 , n17263 , n6364 );
    nor g15161 ( n3541 , n11300 , n29319 );
    or g15162 ( n6856 , n27913 , n23668 );
    xor g15163 ( n22386 , n12053 , n27092 );
    xnor g15164 ( n20526 , n8788 , n22582 );
    not g15165 ( n11833 , n26138 );
    not g15166 ( n3366 , n26024 );
    xnor g15167 ( n30873 , n31794 , n2506 );
    or g15168 ( n4481 , n27348 , n2524 );
    not g15169 ( n6620 , n8268 );
    not g15170 ( n7137 , n31690 );
    or g15171 ( n701 , n2610 , n642 );
    or g15172 ( n20540 , n16255 , n23774 );
    or g15173 ( n4984 , n21996 , n21938 );
    xnor g15174 ( n2424 , n22401 , n14932 );
    and g15175 ( n1075 , n4053 , n9896 );
    xnor g15176 ( n16824 , n29959 , n14788 );
    not g15177 ( n8870 , n3863 );
    xnor g15178 ( n21689 , n31604 , n4213 );
    not g15179 ( n22753 , n25761 );
    xnor g15180 ( n25695 , n12842 , n4453 );
    or g15181 ( n14710 , n16242 , n4998 );
    or g15182 ( n29058 , n15598 , n30658 );
    xnor g15183 ( n1681 , n29477 , n18267 );
    xor g15184 ( n3600 , n27787 , n25275 );
    xnor g15185 ( n11137 , n26871 , n26728 );
    xor g15186 ( n13329 , n18503 , n15228 );
    or g15187 ( n6878 , n8261 , n1975 );
    not g15188 ( n7112 , n23857 );
    not g15189 ( n20269 , n23348 );
    xor g15190 ( n31474 , n1864 , n18730 );
    not g15191 ( n18765 , n27152 );
    xnor g15192 ( n11125 , n31944 , n2191 );
    or g15193 ( n14793 , n11478 , n12684 );
    and g15194 ( n5373 , n5352 , n14050 );
    not g15195 ( n8228 , n15166 );
    or g15196 ( n12311 , n8446 , n14879 );
    xnor g15197 ( n7761 , n3204 , n27689 );
    or g15198 ( n8935 , n16549 , n7717 );
    and g15199 ( n24062 , n898 , n7002 );
    or g15200 ( n22222 , n18120 , n25779 );
    and g15201 ( n22952 , n9599 , n16440 );
    xnor g15202 ( n4891 , n12998 , n22549 );
    xnor g15203 ( n4298 , n1221 , n28006 );
    not g15204 ( n22134 , n3174 );
    not g15205 ( n31748 , n8806 );
    nor g15206 ( n30357 , n28322 , n14518 );
    nor g15207 ( n28094 , n12659 , n4384 );
    xnor g15208 ( n30639 , n4876 , n8335 );
    not g15209 ( n3500 , n13894 );
    not g15210 ( n13864 , n7520 );
    not g15211 ( n12293 , n2934 );
    xnor g15212 ( n16425 , n13723 , n667 );
    and g15213 ( n3950 , n22995 , n24580 );
    xnor g15214 ( n11755 , n15092 , n21474 );
    nor g15215 ( n28542 , n3076 , n9179 );
    or g15216 ( n22034 , n12543 , n6270 );
    or g15217 ( n543 , n5337 , n2369 );
    not g15218 ( n6076 , n28885 );
    nor g15219 ( n237 , n31146 , n8748 );
    xnor g15220 ( n23126 , n4896 , n2556 );
    not g15221 ( n27242 , n14363 );
    xnor g15222 ( n29157 , n7275 , n26430 );
    and g15223 ( n17721 , n18020 , n1090 );
    or g15224 ( n8527 , n14605 , n21856 );
    xnor g15225 ( n15848 , n526 , n25842 );
    and g15226 ( n11251 , n20107 , n7651 );
    nor g15227 ( n14970 , n10058 , n3597 );
    xnor g15228 ( n26119 , n30202 , n2407 );
    or g15229 ( n26850 , n16039 , n8175 );
    not g15230 ( n14144 , n24363 );
    xnor g15231 ( n6487 , n20307 , n26051 );
    nor g15232 ( n286 , n8584 , n1575 );
    or g15233 ( n24284 , n8637 , n16769 );
    and g15234 ( n31975 , n31135 , n28060 );
    not g15235 ( n8468 , n15447 );
    xnor g15236 ( n10190 , n19897 , n15759 );
    or g15237 ( n14889 , n14814 , n23161 );
    not g15238 ( n16870 , n12073 );
    not g15239 ( n16790 , n3859 );
    not g15240 ( n28968 , n16019 );
    and g15241 ( n4892 , n12354 , n3385 );
    xnor g15242 ( n26047 , n13830 , n20927 );
    not g15243 ( n30705 , n27483 );
    xnor g15244 ( n19095 , n22108 , n1733 );
    and g15245 ( n19498 , n1531 , n9714 );
    xnor g15246 ( n23957 , n22891 , n11654 );
    xnor g15247 ( n888 , n24332 , n1776 );
    xnor g15248 ( n6669 , n3689 , n11935 );
    xnor g15249 ( n25362 , n21709 , n509 );
    and g15250 ( n23569 , n10359 , n10854 );
    nor g15251 ( n25417 , n28158 , n20600 );
    xnor g15252 ( n25508 , n20303 , n9587 );
    and g15253 ( n13303 , n30810 , n22961 );
    and g15254 ( n22448 , n21916 , n10722 );
    or g15255 ( n12365 , n13047 , n28805 );
    not g15256 ( n23707 , n12277 );
    and g15257 ( n30362 , n17709 , n26211 );
    or g15258 ( n16959 , n24409 , n29793 );
    xnor g15259 ( n27177 , n30939 , n12713 );
    not g15260 ( n12903 , n26633 );
    xnor g15261 ( n28502 , n25017 , n19981 );
    not g15262 ( n20326 , n19137 );
    xnor g15263 ( n7422 , n25917 , n27354 );
    not g15264 ( n20332 , n25947 );
    nor g15265 ( n4667 , n13454 , n29356 );
    xnor g15266 ( n5014 , n10851 , n16309 );
    not g15267 ( n22970 , n595 );
    or g15268 ( n11596 , n1821 , n3920 );
    not g15269 ( n19646 , n31677 );
    or g15270 ( n28459 , n8747 , n24802 );
    nor g15271 ( n29822 , n3141 , n1283 );
    xnor g15272 ( n4423 , n11690 , n8532 );
    not g15273 ( n27785 , n30414 );
    not g15274 ( n22903 , n6579 );
    not g15275 ( n4648 , n1057 );
    or g15276 ( n7207 , n6792 , n8933 );
    not g15277 ( n20988 , n29963 );
    or g15278 ( n15709 , n20759 , n5933 );
    not g15279 ( n21113 , n13818 );
    not g15280 ( n25332 , n17638 );
    not g15281 ( n3759 , n23023 );
    or g15282 ( n27378 , n31700 , n27924 );
    or g15283 ( n29509 , n4226 , n29415 );
    xnor g15284 ( n13079 , n21207 , n28903 );
    not g15285 ( n15579 , n28600 );
    or g15286 ( n28797 , n16400 , n6234 );
    not g15287 ( n6058 , n26974 );
    not g15288 ( n4161 , n26726 );
    not g15289 ( n7933 , n21186 );
    xor g15290 ( n8593 , n28366 , n27011 );
    not g15291 ( n30061 , n20813 );
    and g15292 ( n21144 , n11214 , n26238 );
    and g15293 ( n6296 , n22592 , n4617 );
    xnor g15294 ( n23308 , n154 , n11905 );
    xnor g15295 ( n5414 , n11724 , n19919 );
    not g15296 ( n5695 , n7313 );
    xnor g15297 ( n28591 , n6036 , n5300 );
    not g15298 ( n20035 , n19344 );
    and g15299 ( n13252 , n25667 , n1124 );
    not g15300 ( n18053 , n17584 );
    not g15301 ( n2352 , n1095 );
    or g15302 ( n15405 , n9850 , n3454 );
    xnor g15303 ( n21810 , n30013 , n948 );
    not g15304 ( n16730 , n12052 );
    or g15305 ( n14077 , n14056 , n13128 );
    and g15306 ( n15770 , n3304 , n21958 );
    not g15307 ( n9825 , n6976 );
    not g15308 ( n17634 , n24782 );
    and g15309 ( n25529 , n16126 , n31637 );
    and g15310 ( n13481 , n31114 , n506 );
    and g15311 ( n1824 , n27017 , n21675 );
    not g15312 ( n27308 , n13433 );
    xor g15313 ( n13344 , n21241 , n10820 );
    and g15314 ( n8352 , n10600 , n6527 );
    xnor g15315 ( n12959 , n1387 , n31617 );
    nor g15316 ( n30647 , n20790 , n28911 );
    xnor g15317 ( n18752 , n3539 , n20697 );
    xnor g15318 ( n26103 , n14737 , n20444 );
    not g15319 ( n28811 , n9888 );
    or g15320 ( n25530 , n2610 , n2933 );
    not g15321 ( n22823 , n9619 );
    xnor g15322 ( n2141 , n16577 , n6612 );
    or g15323 ( n20166 , n7276 , n11465 );
    or g15324 ( n21213 , n21493 , n18045 );
    and g15325 ( n26477 , n24621 , n626 );
    and g15326 ( n10489 , n29327 , n11632 );
    and g15327 ( n21601 , n9093 , n5591 );
    or g15328 ( n25124 , n10676 , n16313 );
    or g15329 ( n23239 , n8486 , n9103 );
    not g15330 ( n27500 , n19440 );
    not g15331 ( n22170 , n20137 );
    xnor g15332 ( n28621 , n32025 , n2447 );
    not g15333 ( n15818 , n8503 );
    or g15334 ( n409 , n27844 , n29338 );
    not g15335 ( n9404 , n10002 );
    not g15336 ( n16920 , n27537 );
    not g15337 ( n10933 , n27420 );
    not g15338 ( n16059 , n8253 );
    and g15339 ( n10573 , n1840 , n27126 );
    and g15340 ( n1674 , n18488 , n25085 );
    xnor g15341 ( n18362 , n30871 , n30002 );
    not g15342 ( n23343 , n14925 );
    or g15343 ( n490 , n30953 , n3007 );
    nor g15344 ( n23053 , n24464 , n9047 );
    xnor g15345 ( n29337 , n16608 , n2864 );
    and g15346 ( n20443 , n15332 , n18586 );
    not g15347 ( n13185 , n5610 );
    xnor g15348 ( n20598 , n19569 , n31896 );
    not g15349 ( n12482 , n20943 );
    or g15350 ( n23531 , n31470 , n740 );
    or g15351 ( n23212 , n13238 , n26274 );
    and g15352 ( n23751 , n5466 , n21397 );
    nor g15353 ( n20918 , n8423 , n10655 );
    or g15354 ( n25449 , n30244 , n959 );
    and g15355 ( n5040 , n10392 , n25719 );
    or g15356 ( n9547 , n6967 , n13544 );
    nor g15357 ( n17619 , n11169 , n6424 );
    xnor g15358 ( n15141 , n4489 , n29132 );
    xnor g15359 ( n29564 , n15169 , n3196 );
    xnor g15360 ( n1458 , n29910 , n25372 );
    not g15361 ( n27384 , n25786 );
    and g15362 ( n13645 , n22457 , n10211 );
    and g15363 ( n3082 , n19848 , n6651 );
    or g15364 ( n23093 , n16199 , n3586 );
    nor g15365 ( n30149 , n7359 , n20493 );
    or g15366 ( n3133 , n20252 , n16801 );
    xnor g15367 ( n28399 , n23301 , n9731 );
    buf g15368 ( n15470 , n23870 );
    xnor g15369 ( n13365 , n22101 , n16512 );
    not g15370 ( n12765 , n6129 );
    or g15371 ( n27323 , n13526 , n29400 );
    not g15372 ( n4159 , n4476 );
    or g15373 ( n19281 , n7823 , n26243 );
    not g15374 ( n1910 , n31034 );
    not g15375 ( n16152 , n31270 );
    not g15376 ( n12619 , n18853 );
    and g15377 ( n10234 , n20376 , n7139 );
    or g15378 ( n13019 , n10385 , n2806 );
    not g15379 ( n21231 , n15360 );
    or g15380 ( n8560 , n21534 , n14074 );
    not g15381 ( n10266 , n10928 );
    and g15382 ( n4189 , n6856 , n16971 );
    not g15383 ( n2717 , n30608 );
    or g15384 ( n16817 , n11813 , n9747 );
    not g15385 ( n30633 , n17882 );
    xnor g15386 ( n8852 , n12925 , n7070 );
    and g15387 ( n28680 , n1063 , n20168 );
    not g15388 ( n3422 , n10653 );
    or g15389 ( n13702 , n10673 , n717 );
    not g15390 ( n19924 , n29187 );
    and g15391 ( n21287 , n18492 , n1715 );
    not g15392 ( n30556 , n13829 );
    xnor g15393 ( n30172 , n16878 , n2092 );
    not g15394 ( n7359 , n17585 );
    nor g15395 ( n11296 , n18850 , n31119 );
    not g15396 ( n20374 , n7191 );
    and g15397 ( n24663 , n19075 , n29247 );
    xnor g15398 ( n25753 , n18929 , n17166 );
    or g15399 ( n6845 , n14577 , n11007 );
    not g15400 ( n23338 , n14018 );
    xor g15401 ( n22905 , n31906 , n3765 );
    and g15402 ( n12780 , n4889 , n14873 );
    not g15403 ( n9757 , n11049 );
    not g15404 ( n1219 , n18207 );
    xnor g15405 ( n17190 , n3220 , n14602 );
    not g15406 ( n24173 , n25991 );
    not g15407 ( n4134 , n16330 );
    or g15408 ( n27607 , n5153 , n10464 );
    or g15409 ( n12098 , n13700 , n9699 );
    or g15410 ( n13445 , n13635 , n8120 );
    not g15411 ( n13281 , n8507 );
    or g15412 ( n30350 , n6626 , n3412 );
    or g15413 ( n31207 , n12443 , n15315 );
    xor g15414 ( n2545 , n26537 , n18117 );
    xnor g15415 ( n13470 , n27317 , n14489 );
    xnor g15416 ( n30249 , n10022 , n21649 );
    xnor g15417 ( n31246 , n26050 , n19727 );
    not g15418 ( n1130 , n16934 );
    or g15419 ( n25592 , n14425 , n20164 );
    and g15420 ( n12559 , n19510 , n5936 );
    not g15421 ( n19457 , n7220 );
    not g15422 ( n20489 , n19315 );
    not g15423 ( n21742 , n10790 );
    not g15424 ( n23767 , n16794 );
    xnor g15425 ( n8980 , n6791 , n21527 );
    or g15426 ( n12362 , n9216 , n23111 );
    and g15427 ( n8525 , n15029 , n9479 );
    xnor g15428 ( n16776 , n2257 , n27748 );
    xnor g15429 ( n11756 , n2073 , n26329 );
    and g15430 ( n29674 , n22267 , n11957 );
    or g15431 ( n25942 , n20469 , n21976 );
    not g15432 ( n2292 , n8862 );
    not g15433 ( n17044 , n31115 );
    xnor g15434 ( n13417 , n14505 , n9215 );
    xnor g15435 ( n1887 , n10807 , n27302 );
    nor g15436 ( n3032 , n22019 , n850 );
    nor g15437 ( n10594 , n13454 , n4499 );
    and g15438 ( n11406 , n14132 , n24525 );
    or g15439 ( n30835 , n14764 , n9201 );
    and g15440 ( n3371 , n985 , n21876 );
    not g15441 ( n11094 , n2862 );
    or g15442 ( n24156 , n22608 , n23201 );
    and g15443 ( n22397 , n2612 , n3594 );
    and g15444 ( n31044 , n24200 , n10654 );
    nor g15445 ( n10276 , n18800 , n17863 );
    or g15446 ( n2293 , n4844 , n4009 );
    not g15447 ( n31038 , n14809 );
    or g15448 ( n31508 , n11711 , n25033 );
    or g15449 ( n12705 , n994 , n5068 );
    xnor g15450 ( n31494 , n28234 , n17851 );
    or g15451 ( n24189 , n12860 , n28712 );
    xnor g15452 ( n26150 , n24762 , n9939 );
    or g15453 ( n20264 , n21043 , n16964 );
    not g15454 ( n13203 , n28507 );
    or g15455 ( n609 , n28096 , n989 );
    nor g15456 ( n19190 , n13700 , n12802 );
    xnor g15457 ( n22469 , n3225 , n1285 );
    not g15458 ( n18707 , n4995 );
    nor g15459 ( n27943 , n16132 , n13817 );
    or g15460 ( n13884 , n17913 , n15792 );
    or g15461 ( n13709 , n14287 , n30575 );
    not g15462 ( n6819 , n23035 );
    not g15463 ( n1267 , n17265 );
    xnor g15464 ( n695 , n27061 , n16166 );
    not g15465 ( n28114 , n3068 );
    or g15466 ( n20076 , n25625 , n30981 );
    xnor g15467 ( n22243 , n632 , n4257 );
    xnor g15468 ( n10612 , n30022 , n29668 );
    xnor g15469 ( n31015 , n19019 , n25199 );
    xor g15470 ( n13495 , n7805 , n28891 );
    xnor g15471 ( n28019 , n20687 , n17086 );
    not g15472 ( n23667 , n8713 );
    xnor g15473 ( n5227 , n17664 , n30373 );
    and g15474 ( n15516 , n9028 , n24601 );
    not g15475 ( n21609 , n1484 );
    or g15476 ( n23600 , n30685 , n15849 );
    xnor g15477 ( n23635 , n138 , n3297 );
    or g15478 ( n23190 , n25943 , n11210 );
    or g15479 ( n9666 , n7027 , n4837 );
    not g15480 ( n12897 , n31875 );
    nor g15481 ( n1899 , n11302 , n6955 );
    nor g15482 ( n24579 , n31365 , n21579 );
    or g15483 ( n2769 , n21344 , n25418 );
    or g15484 ( n6691 , n5161 , n12811 );
    and g15485 ( n25484 , n25584 , n2305 );
    nor g15486 ( n31357 , n594 , n9537 );
    xnor g15487 ( n8762 , n22522 , n2001 );
    not g15488 ( n15836 , n8906 );
    not g15489 ( n2815 , n15479 );
    xnor g15490 ( n30667 , n24826 , n13549 );
    or g15491 ( n5849 , n28656 , n23610 );
    nor g15492 ( n4550 , n1537 , n21610 );
    not g15493 ( n19974 , n5114 );
    not g15494 ( n12418 , n6260 );
    and g15495 ( n12510 , n6829 , n15375 );
    not g15496 ( n15674 , n23082 );
    xnor g15497 ( n31083 , n10111 , n4402 );
    not g15498 ( n2562 , n1585 );
    or g15499 ( n21825 , n2432 , n3759 );
    nor g15500 ( n22146 , n27077 , n7496 );
    xnor g15501 ( n12584 , n29764 , n29604 );
    and g15502 ( n12278 , n15331 , n18383 );
    not g15503 ( n13739 , n3170 );
    nor g15504 ( n3015 , n3634 , n19618 );
    not g15505 ( n2018 , n8680 );
    xnor g15506 ( n15164 , n15959 , n25557 );
    nor g15507 ( n29599 , n19254 , n13188 );
    xnor g15508 ( n30897 , n15186 , n22522 );
    and g15509 ( n30668 , n17742 , n5631 );
    nor g15510 ( n21640 , n27498 , n23889 );
    xnor g15511 ( n21174 , n23617 , n14471 );
    xnor g15512 ( n18925 , n25855 , n2300 );
    not g15513 ( n20115 , n29236 );
    and g15514 ( n18343 , n4017 , n21103 );
    and g15515 ( n1502 , n16993 , n10116 );
    xnor g15516 ( n14627 , n18633 , n24345 );
    xnor g15517 ( n26376 , n1287 , n25047 );
    or g15518 ( n5393 , n25482 , n6484 );
    xnor g15519 ( n1202 , n910 , n19658 );
    not g15520 ( n23579 , n24662 );
    or g15521 ( n27692 , n10114 , n7934 );
    xnor g15522 ( n18107 , n12958 , n9388 );
    or g15523 ( n29429 , n29503 , n29689 );
    or g15524 ( n16896 , n26654 , n3100 );
    nor g15525 ( n2643 , n14520 , n28281 );
    and g15526 ( n18492 , n13590 , n1640 );
    and g15527 ( n12808 , n24109 , n28969 );
    and g15528 ( n13713 , n13623 , n29858 );
    not g15529 ( n18316 , n327 );
    and g15530 ( n23581 , n2200 , n29294 );
    not g15531 ( n13948 , n26894 );
    xnor g15532 ( n20753 , n5961 , n19769 );
    or g15533 ( n15764 , n24924 , n17117 );
    not g15534 ( n5190 , n26185 );
    and g15535 ( n29915 , n15428 , n18513 );
    or g15536 ( n25537 , n803 , n30635 );
    and g15537 ( n23544 , n17503 , n22976 );
    or g15538 ( n6272 , n25147 , n2297 );
    xnor g15539 ( n3423 , n12933 , n9118 );
    xnor g15540 ( n1722 , n20053 , n29269 );
    or g15541 ( n22741 , n4789 , n27089 );
    or g15542 ( n24378 , n1566 , n26562 );
    not g15543 ( n18764 , n8321 );
    not g15544 ( n30208 , n12765 );
    not g15545 ( n14333 , n7621 );
    and g15546 ( n11917 , n30217 , n5947 );
    and g15547 ( n9907 , n13696 , n30049 );
    or g15548 ( n20851 , n1195 , n3163 );
    and g15549 ( n13119 , n19639 , n16394 );
    and g15550 ( n30568 , n7063 , n10397 );
    not g15551 ( n30858 , n23701 );
    not g15552 ( n3090 , n26731 );
    and g15553 ( n17178 , n19045 , n24508 );
    or g15554 ( n12826 , n30716 , n7893 );
    not g15555 ( n3160 , n14239 );
    xor g15556 ( n7697 , n19111 , n17015 );
    xnor g15557 ( n9908 , n11844 , n1280 );
    or g15558 ( n17047 , n26326 , n27659 );
    or g15559 ( n27369 , n29462 , n23472 );
    not g15560 ( n14705 , n26451 );
    xnor g15561 ( n30811 , n14992 , n23561 );
    and g15562 ( n29152 , n10362 , n14672 );
    nor g15563 ( n18953 , n15577 , n27966 );
    or g15564 ( n30545 , n14789 , n5240 );
    and g15565 ( n3007 , n17237 , n22105 );
    or g15566 ( n23278 , n664 , n6962 );
    or g15567 ( n2168 , n18464 , n31435 );
    not g15568 ( n28350 , n622 );
    xnor g15569 ( n2950 , n29776 , n23414 );
    xnor g15570 ( n19858 , n19728 , n14503 );
    xnor g15571 ( n8563 , n31971 , n6645 );
    xnor g15572 ( n11555 , n24220 , n7479 );
    xnor g15573 ( n13372 , n4761 , n17731 );
    not g15574 ( n9233 , n30065 );
    not g15575 ( n7929 , n16870 );
    and g15576 ( n27618 , n12979 , n2870 );
    xnor g15577 ( n3156 , n2758 , n9037 );
    xnor g15578 ( n30940 , n16851 , n13980 );
    nor g15579 ( n11892 , n2628 , n17209 );
    xnor g15580 ( n29101 , n15731 , n7380 );
    xnor g15581 ( n13583 , n2522 , n23611 );
    not g15582 ( n17210 , n20943 );
    or g15583 ( n31268 , n6071 , n13571 );
    xnor g15584 ( n23804 , n22579 , n9342 );
    or g15585 ( n29018 , n22060 , n18125 );
    and g15586 ( n16064 , n28561 , n7016 );
    xnor g15587 ( n29180 , n15376 , n9398 );
    and g15588 ( n19128 , n13098 , n24516 );
    and g15589 ( n16941 , n19784 , n11707 );
    or g15590 ( n23033 , n15102 , n7917 );
    not g15591 ( n27503 , n21265 );
    buf g15592 ( n8360 , n11206 );
    xnor g15593 ( n6577 , n7687 , n30268 );
    or g15594 ( n3476 , n15767 , n26784 );
    or g15595 ( n28253 , n15296 , n22299 );
    xnor g15596 ( n29351 , n2619 , n24448 );
    and g15597 ( n4378 , n22321 , n20173 );
    not g15598 ( n19120 , n6043 );
    not g15599 ( n27559 , n23083 );
    or g15600 ( n29446 , n18602 , n18790 );
    not g15601 ( n20380 , n22641 );
    or g15602 ( n25119 , n3757 , n9444 );
    or g15603 ( n9229 , n20760 , n30565 );
    and g15604 ( n15004 , n28470 , n31889 );
    or g15605 ( n9947 , n9141 , n2815 );
    nor g15606 ( n18219 , n12312 , n10737 );
    buf g15607 ( n10841 , n14102 );
    not g15608 ( n16342 , n3688 );
    or g15609 ( n15001 , n1478 , n22370 );
    and g15610 ( n5476 , n7524 , n2302 );
    xnor g15611 ( n15787 , n13386 , n26593 );
    not g15612 ( n26085 , n10899 );
    not g15613 ( n29166 , n14155 );
    xnor g15614 ( n10064 , n2596 , n9948 );
    nor g15615 ( n139 , n20311 , n17652 );
    nor g15616 ( n20095 , n7434 , n3106 );
    xnor g15617 ( n27237 , n25648 , n17007 );
    and g15618 ( n8022 , n2229 , n5186 );
    xnor g15619 ( n24466 , n18835 , n1213 );
    xnor g15620 ( n21412 , n26696 , n8505 );
    or g15621 ( n3598 , n28100 , n12633 );
    not g15622 ( n11908 , n11788 );
    not g15623 ( n15479 , n8117 );
    or g15624 ( n13368 , n21881 , n32016 );
    not g15625 ( n21564 , n21003 );
    not g15626 ( n28288 , n29991 );
    nor g15627 ( n27335 , n18996 , n9548 );
    and g15628 ( n25800 , n24105 , n24432 );
    or g15629 ( n16889 , n11867 , n25896 );
    not g15630 ( n11482 , n11639 );
    and g15631 ( n16231 , n14354 , n21933 );
    not g15632 ( n5209 , n12105 );
    xnor g15633 ( n24866 , n8806 , n15222 );
    not g15634 ( n18996 , n8426 );
    nor g15635 ( n15366 , n10202 , n3436 );
    not g15636 ( n24313 , n3498 );
    and g15637 ( n7695 , n611 , n20362 );
    not g15638 ( n10394 , n22405 );
    xnor g15639 ( n4547 , n16887 , n14112 );
    or g15640 ( n29610 , n13329 , n16660 );
    and g15641 ( n22189 , n9921 , n9384 );
    not g15642 ( n6010 , n28164 );
    not g15643 ( n30242 , n27005 );
    nor g15644 ( n24983 , n28391 , n1647 );
    xor g15645 ( n22065 , n5772 , n26918 );
    not g15646 ( n2533 , n14318 );
    not g15647 ( n1812 , n22308 );
    or g15648 ( n20221 , n31446 , n10294 );
    or g15649 ( n12476 , n27560 , n2890 );
    xnor g15650 ( n26392 , n30831 , n24794 );
    nor g15651 ( n19412 , n24111 , n4144 );
    xnor g15652 ( n17172 , n16375 , n16674 );
    or g15653 ( n668 , n22099 , n22890 );
    not g15654 ( n30200 , n29343 );
    and g15655 ( n2874 , n25309 , n15882 );
    xnor g15656 ( n6977 , n4155 , n15094 );
    or g15657 ( n13294 , n9934 , n29546 );
    xnor g15658 ( n15617 , n20638 , n27248 );
    xnor g15659 ( n12576 , n5783 , n10393 );
    nor g15660 ( n14850 , n6123 , n1590 );
    not g15661 ( n27093 , n7722 );
    or g15662 ( n1662 , n28939 , n19927 );
    xnor g15663 ( n26547 , n20136 , n22813 );
    or g15664 ( n24379 , n9729 , n31080 );
    nor g15665 ( n9695 , n26066 , n4602 );
    and g15666 ( n11936 , n22061 , n24677 );
    xnor g15667 ( n11063 , n879 , n7871 );
    xnor g15668 ( n23605 , n29380 , n28433 );
    not g15669 ( n23713 , n24896 );
    xnor g15670 ( n31723 , n23618 , n20472 );
    xnor g15671 ( n25431 , n23580 , n31037 );
    and g15672 ( n9974 , n24809 , n6025 );
    xnor g15673 ( n17822 , n29237 , n6534 );
    and g15674 ( n3718 , n28042 , n17817 );
    or g15675 ( n12927 , n14944 , n21915 );
    xnor g15676 ( n3622 , n20041 , n757 );
    xnor g15677 ( n31824 , n24140 , n5666 );
    not g15678 ( n4599 , n10146 );
    xnor g15679 ( n4482 , n10512 , n2242 );
    or g15680 ( n21427 , n12568 , n9615 );
    and g15681 ( n7048 , n29607 , n28709 );
    or g15682 ( n9046 , n10605 , n17603 );
    not g15683 ( n9915 , n19425 );
    not g15684 ( n8346 , n24598 );
    and g15685 ( n15667 , n3638 , n9033 );
    and g15686 ( n31768 , n200 , n5693 );
    or g15687 ( n21117 , n561 , n26555 );
    and g15688 ( n19123 , n22289 , n16878 );
    not g15689 ( n14282 , n3752 );
    xnor g15690 ( n3455 , n13714 , n2177 );
    not g15691 ( n8139 , n16498 );
    not g15692 ( n6188 , n995 );
    and g15693 ( n23034 , n24924 , n17117 );
    and g15694 ( n30966 , n8055 , n27631 );
    not g15695 ( n5202 , n14425 );
    not g15696 ( n23252 , n13330 );
    and g15697 ( n30780 , n7474 , n22414 );
    not g15698 ( n20971 , n13640 );
    xnor g15699 ( n9159 , n27900 , n25295 );
    xnor g15700 ( n25788 , n8714 , n13526 );
    not g15701 ( n3081 , n26067 );
    xnor g15702 ( n12807 , n31078 , n30201 );
    or g15703 ( n4787 , n25939 , n15518 );
    or g15704 ( n29653 , n27049 , n7807 );
    xnor g15705 ( n8566 , n11143 , n1247 );
    not g15706 ( n9642 , n6686 );
    nor g15707 ( n29198 , n19069 , n22606 );
    and g15708 ( n8842 , n24706 , n28251 );
    not g15709 ( n2674 , n8256 );
    not g15710 ( n18609 , n24201 );
    not g15711 ( n27746 , n4159 );
    or g15712 ( n13832 , n19870 , n18109 );
    and g15713 ( n8812 , n29410 , n19278 );
    xnor g15714 ( n12077 , n6471 , n31882 );
    nor g15715 ( n11268 , n19282 , n31496 );
    not g15716 ( n22440 , n4052 );
    nor g15717 ( n4566 , n12941 , n26687 );
    nor g15718 ( n2138 , n28252 , n16273 );
    or g15719 ( n896 , n5490 , n12102 );
    or g15720 ( n2441 , n5395 , n10930 );
    or g15721 ( n30072 , n27885 , n8576 );
    and g15722 ( n789 , n3886 , n26093 );
    and g15723 ( n6576 , n1297 , n20527 );
    and g15724 ( n25644 , n4926 , n26929 );
    xor g15725 ( n12263 , n14185 , n3863 );
    not g15726 ( n20421 , n24802 );
    or g15727 ( n5210 , n29526 , n16796 );
    and g15728 ( n30745 , n19787 , n30694 );
    not g15729 ( n27646 , n20014 );
    xnor g15730 ( n9985 , n25767 , n31263 );
    not g15731 ( n530 , n21707 );
    xnor g15732 ( n5983 , n16889 , n6595 );
    xnor g15733 ( n5046 , n21493 , n7009 );
    and g15734 ( n6749 , n15959 , n23506 );
    and g15735 ( n9293 , n11431 , n16634 );
    not g15736 ( n7325 , n847 );
    xor g15737 ( n1591 , n17738 , n9733 );
    not g15738 ( n4715 , n25447 );
    and g15739 ( n27388 , n21477 , n8721 );
    not g15740 ( n1444 , n18516 );
    xnor g15741 ( n23653 , n22047 , n16930 );
    xnor g15742 ( n31264 , n22955 , n22730 );
    xnor g15743 ( n27737 , n1536 , n1742 );
    xnor g15744 ( n31370 , n22252 , n26229 );
    or g15745 ( n15355 , n18265 , n20052 );
    not g15746 ( n30148 , n15745 );
    not g15747 ( n7218 , n13494 );
    and g15748 ( n24751 , n13217 , n20272 );
    and g15749 ( n23951 , n29146 , n11090 );
    and g15750 ( n1163 , n1490 , n8368 );
    or g15751 ( n6413 , n3696 , n16842 );
    xnor g15752 ( n16070 , n9755 , n11811 );
    and g15753 ( n6542 , n20950 , n7914 );
    or g15754 ( n18601 , n3620 , n5814 );
    xnor g15755 ( n8180 , n7121 , n12077 );
    xnor g15756 ( n31811 , n3763 , n20630 );
    xnor g15757 ( n5416 , n12522 , n24569 );
    or g15758 ( n29577 , n3134 , n4329 );
    not g15759 ( n13005 , n20146 );
    and g15760 ( n29000 , n12115 , n26041 );
    not g15761 ( n453 , n3085 );
    nor g15762 ( n14183 , n27883 , n26460 );
    xnor g15763 ( n5820 , n26688 , n17864 );
    xnor g15764 ( n26228 , n8122 , n15083 );
    xnor g15765 ( n6334 , n96 , n5757 );
    xnor g15766 ( n12933 , n7597 , n12224 );
    nor g15767 ( n7401 , n1518 , n10676 );
    xnor g15768 ( n20320 , n11764 , n2301 );
    or g15769 ( n11429 , n14830 , n8084 );
    or g15770 ( n2672 , n17973 , n14006 );
    not g15771 ( n18506 , n22512 );
    and g15772 ( n13248 , n5740 , n7954 );
    not g15773 ( n19700 , n996 );
    and g15774 ( n20946 , n6694 , n10826 );
    or g15775 ( n22791 , n31240 , n29651 );
    nor g15776 ( n9496 , n2694 , n8939 );
    and g15777 ( n17523 , n23115 , n24837 );
    and g15778 ( n24832 , n25792 , n27638 );
    and g15779 ( n12003 , n9364 , n13783 );
    or g15780 ( n27047 , n2715 , n20255 );
    xnor g15781 ( n9449 , n27452 , n11729 );
    or g15782 ( n23560 , n20751 , n27203 );
    not g15783 ( n16991 , n11187 );
    or g15784 ( n30638 , n4574 , n18102 );
    nor g15785 ( n16467 , n14796 , n12284 );
    not g15786 ( n16617 , n12684 );
    not g15787 ( n9 , n1073 );
    or g15788 ( n21864 , n27897 , n12544 );
    xnor g15789 ( n391 , n31382 , n10151 );
    or g15790 ( n7976 , n18595 , n2937 );
    xnor g15791 ( n27141 , n1805 , n29646 );
    xnor g15792 ( n28040 , n17177 , n16881 );
    xnor g15793 ( n21475 , n30887 , n28983 );
    and g15794 ( n9887 , n10298 , n25232 );
    not g15795 ( n5501 , n7458 );
    not g15796 ( n6968 , n27272 );
    and g15797 ( n11294 , n27740 , n31885 );
    not g15798 ( n20625 , n23620 );
    xnor g15799 ( n11039 , n26719 , n28451 );
    or g15800 ( n23794 , n9791 , n20951 );
    not g15801 ( n2000 , n30746 );
    nor g15802 ( n13412 , n12207 , n14738 );
    and g15803 ( n26717 , n6805 , n17359 );
    xnor g15804 ( n4344 , n3246 , n31198 );
    and g15805 ( n195 , n25664 , n21939 );
    not g15806 ( n20600 , n8014 );
    xnor g15807 ( n21790 , n6030 , n21332 );
    nor g15808 ( n13411 , n30201 , n12175 );
    xnor g15809 ( n28754 , n26372 , n21703 );
    or g15810 ( n17858 , n13591 , n19877 );
    or g15811 ( n27614 , n30038 , n17178 );
    or g15812 ( n28905 , n18815 , n430 );
    xnor g15813 ( n12275 , n29618 , n1771 );
    nor g15814 ( n14814 , n16200 , n16342 );
    xnor g15815 ( n11370 , n10066 , n20487 );
    not g15816 ( n21522 , n13640 );
    xnor g15817 ( n2190 , n14853 , n22851 );
    xnor g15818 ( n8344 , n9853 , n2704 );
    xnor g15819 ( n14118 , n18288 , n28712 );
    not g15820 ( n20371 , n26261 );
    or g15821 ( n23816 , n5019 , n394 );
    not g15822 ( n12279 , n14201 );
    or g15823 ( n8837 , n10208 , n14270 );
    nor g15824 ( n30680 , n19372 , n10664 );
    xnor g15825 ( n4267 , n21731 , n4466 );
    not g15826 ( n9353 , n2782 );
    and g15827 ( n29240 , n18964 , n23537 );
    not g15828 ( n2044 , n12024 );
    and g15829 ( n1902 , n9276 , n29974 );
    not g15830 ( n31051 , n15807 );
    or g15831 ( n10648 , n21918 , n6651 );
    or g15832 ( n11135 , n23455 , n18065 );
    or g15833 ( n21666 , n14624 , n11973 );
    and g15834 ( n5042 , n27854 , n13834 );
    or g15835 ( n10035 , n19545 , n11237 );
    or g15836 ( n25271 , n31586 , n15862 );
    xnor g15837 ( n9837 , n29082 , n13688 );
    not g15838 ( n4012 , n30633 );
    not g15839 ( n19558 , n4128 );
    or g15840 ( n20077 , n5750 , n25824 );
    and g15841 ( n26925 , n333 , n1074 );
    and g15842 ( n31719 , n11976 , n1869 );
    and g15843 ( n5571 , n9665 , n24462 );
    not g15844 ( n29064 , n24104 );
    not g15845 ( n9241 , n30044 );
    xnor g15846 ( n17318 , n11900 , n16083 );
    xnor g15847 ( n14507 , n4455 , n13440 );
    not g15848 ( n18983 , n17026 );
    or g15849 ( n4337 , n19466 , n504 );
    nor g15850 ( n15992 , n2301 , n25093 );
    not g15851 ( n19082 , n7433 );
    xnor g15852 ( n29745 , n1641 , n26159 );
    and g15853 ( n6459 , n8071 , n22736 );
    not g15854 ( n19087 , n12790 );
    or g15855 ( n23895 , n16032 , n7585 );
    and g15856 ( n19690 , n23392 , n23929 );
    or g15857 ( n4217 , n4832 , n14923 );
    not g15858 ( n4864 , n7342 );
    not g15859 ( n1942 , n3485 );
    not g15860 ( n28147 , n24281 );
    nor g15861 ( n16556 , n23899 , n27057 );
    xnor g15862 ( n25509 , n13943 , n28541 );
    not g15863 ( n13259 , n9118 );
    not g15864 ( n7547 , n26410 );
    xor g15865 ( n19137 , n17411 , n22678 );
    xnor g15866 ( n11 , n27791 , n22348 );
    or g15867 ( n9100 , n3822 , n5822 );
    or g15868 ( n23477 , n24350 , n11290 );
    xnor g15869 ( n4733 , n491 , n5967 );
    or g15870 ( n11432 , n16645 , n744 );
    xnor g15871 ( n5840 , n14770 , n21767 );
    nor g15872 ( n14211 , n4676 , n8396 );
    nor g15873 ( n4732 , n20667 , n25299 );
    not g15874 ( n11933 , n9862 );
    not g15875 ( n6619 , n27207 );
    not g15876 ( n204 , n20058 );
    xnor g15877 ( n31048 , n19887 , n11597 );
    or g15878 ( n31946 , n2100 , n6118 );
    xnor g15879 ( n1618 , n29825 , n24074 );
    not g15880 ( n18157 , n11218 );
    or g15881 ( n11558 , n24383 , n21710 );
    xnor g15882 ( n20929 , n18864 , n13291 );
    xnor g15883 ( n20917 , n12705 , n15544 );
    not g15884 ( n18378 , n7315 );
    or g15885 ( n21788 , n10105 , n9549 );
    or g15886 ( n25126 , n21206 , n29487 );
    and g15887 ( n17699 , n1552 , n14954 );
    or g15888 ( n4314 , n24396 , n591 );
    xnor g15889 ( n20555 , n20357 , n7720 );
    not g15890 ( n25499 , n21454 );
    not g15891 ( n15017 , n12542 );
    and g15892 ( n12840 , n10533 , n26440 );
    not g15893 ( n6210 , n15664 );
    and g15894 ( n30520 , n27822 , n22613 );
    not g15895 ( n28444 , n19558 );
    xnor g15896 ( n13073 , n21974 , n24147 );
    not g15897 ( n21091 , n16130 );
    not g15898 ( n26686 , n23218 );
    nor g15899 ( n31780 , n13471 , n29046 );
    or g15900 ( n15167 , n1269 , n10920 );
    xnor g15901 ( n21632 , n23672 , n3400 );
    xnor g15902 ( n20501 , n5388 , n1856 );
    xnor g15903 ( n28169 , n11492 , n13244 );
    not g15904 ( n16302 , n13854 );
    or g15905 ( n11376 , n8714 , n675 );
    and g15906 ( n25315 , n7234 , n23223 );
    and g15907 ( n12738 , n7306 , n25249 );
    or g15908 ( n9622 , n664 , n11050 );
    or g15909 ( n20036 , n20552 , n11434 );
    not g15910 ( n25387 , n13568 );
    nor g15911 ( n19955 , n21310 , n10210 );
    xor g15912 ( n31503 , n440 , n23308 );
    or g15913 ( n3644 , n19871 , n29661 );
    not g15914 ( n28546 , n22233 );
    xnor g15915 ( n21313 , n27611 , n28890 );
    xnor g15916 ( n2605 , n11894 , n9146 );
    xnor g15917 ( n9709 , n24149 , n23052 );
    or g15918 ( n17581 , n17274 , n7260 );
    nor g15919 ( n18008 , n28509 , n18161 );
    or g15920 ( n27422 , n24412 , n24099 );
    and g15921 ( n7528 , n6359 , n20846 );
    not g15922 ( n17906 , n15365 );
    xor g15923 ( n6465 , n30137 , n2764 );
    or g15924 ( n6747 , n30602 , n3375 );
    and g15925 ( n119 , n103 , n23935 );
    or g15926 ( n13869 , n21584 , n13130 );
    or g15927 ( n24357 , n18415 , n321 );
    xnor g15928 ( n24841 , n22950 , n7903 );
    xor g15929 ( n8017 , n28073 , n11886 );
    and g15930 ( n7966 , n28082 , n25875 );
    xnor g15931 ( n8944 , n31768 , n13981 );
    or g15932 ( n27485 , n3090 , n8845 );
    not g15933 ( n17173 , n4568 );
    xnor g15934 ( n17540 , n29056 , n3197 );
    not g15935 ( n2041 , n17880 );
    xnor g15936 ( n5275 , n8587 , n6498 );
    xnor g15937 ( n16729 , n26107 , n13257 );
    or g15938 ( n26990 , n3887 , n4018 );
    xnor g15939 ( n16156 , n3810 , n10433 );
    xnor g15940 ( n8145 , n28139 , n5754 );
    nor g15941 ( n1264 , n23334 , n23680 );
    nor g15942 ( n10268 , n9424 , n29323 );
    nor g15943 ( n2050 , n19615 , n16406 );
    and g15944 ( n7873 , n13007 , n16165 );
    or g15945 ( n3617 , n12803 , n5746 );
    nor g15946 ( n8768 , n23419 , n13376 );
    or g15947 ( n21791 , n17206 , n30191 );
    not g15948 ( n24489 , n20798 );
    not g15949 ( n23528 , n18418 );
    not g15950 ( n30607 , n28402 );
    or g15951 ( n6344 , n30688 , n1073 );
    nor g15952 ( n14172 , n5561 , n28914 );
    not g15953 ( n10944 , n22573 );
    buf g15954 ( n15669 , n31337 );
    or g15955 ( n28015 , n14313 , n20464 );
    xnor g15956 ( n30363 , n13061 , n16583 );
    nor g15957 ( n7171 , n4054 , n7214 );
    or g15958 ( n2873 , n12070 , n4040 );
    xnor g15959 ( n7133 , n16811 , n25364 );
    or g15960 ( n20559 , n24008 , n27914 );
    not g15961 ( n4144 , n14102 );
    not g15962 ( n17487 , n5949 );
    xnor g15963 ( n8460 , n17984 , n9568 );
    xnor g15964 ( n27708 , n21575 , n20092 );
    xnor g15965 ( n18803 , n7738 , n20782 );
    xnor g15966 ( n25665 , n1473 , n19581 );
    nor g15967 ( n10376 , n29715 , n5274 );
    or g15968 ( n29913 , n19211 , n11928 );
    and g15969 ( n709 , n8999 , n15604 );
    xor g15970 ( n5306 , n22308 , n12034 );
    xnor g15971 ( n26908 , n22312 , n7671 );
    or g15972 ( n18896 , n11927 , n18643 );
    or g15973 ( n29396 , n18371 , n6685 );
    xnor g15974 ( n20129 , n14623 , n27546 );
    not g15975 ( n27021 , n20106 );
    not g15976 ( n20608 , n4358 );
    not g15977 ( n6030 , n13103 );
    and g15978 ( n27140 , n23553 , n882 );
    nor g15979 ( n20499 , n29876 , n29940 );
    xnor g15980 ( n25884 , n13026 , n21409 );
    and g15981 ( n24642 , n17247 , n18680 );
    nor g15982 ( n17732 , n5631 , n28106 );
    or g15983 ( n18911 , n24038 , n15682 );
    and g15984 ( n702 , n2365 , n13045 );
    not g15985 ( n20463 , n30245 );
    and g15986 ( n2886 , n26582 , n29809 );
    xnor g15987 ( n2558 , n8492 , n6988 );
    xnor g15988 ( n922 , n13319 , n21464 );
    or g15989 ( n19900 , n21473 , n25829 );
    and g15990 ( n17467 , n25900 , n11771 );
    or g15991 ( n21108 , n19495 , n14224 );
    not g15992 ( n26884 , n7564 );
    and g15993 ( n22810 , n2625 , n11007 );
    nor g15994 ( n5488 , n18002 , n31897 );
    not g15995 ( n6078 , n20820 );
    or g15996 ( n22923 , n2576 , n10916 );
    not g15997 ( n15967 , n24271 );
    not g15998 ( n27684 , n27737 );
    xnor g15999 ( n412 , n28983 , n8584 );
    or g16000 ( n2633 , n28249 , n15440 );
    not g16001 ( n10564 , n17151 );
    and g16002 ( n15552 , n26140 , n12285 );
    xnor g16003 ( n12441 , n27197 , n28472 );
    not g16004 ( n4318 , n8909 );
    and g16005 ( n19019 , n26881 , n27905 );
    not g16006 ( n27651 , n17548 );
    not g16007 ( n18349 , n11354 );
    not g16008 ( n28837 , n14712 );
    xnor g16009 ( n8902 , n4867 , n26492 );
    xor g16010 ( n9769 , n18874 , n18536 );
    not g16011 ( n11517 , n1346 );
    or g16012 ( n10 , n30676 , n4728 );
    or g16013 ( n8795 , n22122 , n4256 );
    or g16014 ( n18233 , n26976 , n8391 );
    or g16015 ( n13881 , n29152 , n507 );
    and g16016 ( n11443 , n9741 , n6239 );
    and g16017 ( n21797 , n4373 , n10132 );
    xnor g16018 ( n9775 , n24621 , n626 );
    not g16019 ( n16779 , n6874 );
    not g16020 ( n14318 , n11447 );
    and g16021 ( n16954 , n21199 , n7003 );
    and g16022 ( n24012 , n16175 , n3382 );
    not g16023 ( n17778 , n10218 );
    not g16024 ( n29529 , n17692 );
    not g16025 ( n5479 , n158 );
    nor g16026 ( n9765 , n28111 , n17624 );
    xnor g16027 ( n21013 , n29664 , n12768 );
    xnor g16028 ( n17033 , n14795 , n22866 );
    not g16029 ( n4690 , n1783 );
    xnor g16030 ( n4051 , n26782 , n17734 );
    or g16031 ( n20145 , n14033 , n6823 );
    not g16032 ( n31465 , n3949 );
    or g16033 ( n30354 , n25004 , n18986 );
    xnor g16034 ( n24622 , n28549 , n23567 );
    not g16035 ( n25174 , n5882 );
    buf g16036 ( n19790 , n19056 );
    xnor g16037 ( n19108 , n9184 , n5148 );
    not g16038 ( n12353 , n15865 );
    and g16039 ( n20405 , n7886 , n7207 );
    xnor g16040 ( n9885 , n19806 , n18094 );
    and g16041 ( n31302 , n15928 , n22107 );
    not g16042 ( n26354 , n30121 );
    or g16043 ( n27631 , n16558 , n10334 );
    and g16044 ( n4125 , n13225 , n16386 );
    and g16045 ( n25855 , n13139 , n5978 );
    and g16046 ( n24884 , n31729 , n11581 );
    not g16047 ( n20294 , n9354 );
    xnor g16048 ( n1686 , n30326 , n9414 );
    xnor g16049 ( n27895 , n9668 , n28854 );
    and g16050 ( n15251 , n12775 , n7042 );
    nor g16051 ( n14150 , n2543 , n5974 );
    xnor g16052 ( n1944 , n31568 , n30238 );
    not g16053 ( n31800 , n9788 );
    xnor g16054 ( n7308 , n24019 , n6145 );
    not g16055 ( n10214 , n17688 );
    or g16056 ( n22032 , n16565 , n29413 );
    not g16057 ( n23051 , n5432 );
    or g16058 ( n29511 , n5268 , n924 );
    xnor g16059 ( n18980 , n16501 , n5592 );
    or g16060 ( n5087 , n20489 , n13060 );
    or g16061 ( n26104 , n29040 , n12003 );
    xnor g16062 ( n22389 , n1177 , n31470 );
    and g16063 ( n8059 , n6323 , n3827 );
    or g16064 ( n7737 , n4058 , n18610 );
    not g16065 ( n16890 , n125 );
    not g16066 ( n30717 , n6254 );
    nor g16067 ( n23590 , n9318 , n8919 );
    not g16068 ( n18700 , n22022 );
    not g16069 ( n19071 , n27770 );
    not g16070 ( n5594 , n25527 );
    not g16071 ( n17037 , n3307 );
    not g16072 ( n25290 , n8986 );
    not g16073 ( n12801 , n20021 );
    and g16074 ( n8215 , n16337 , n12088 );
    not g16075 ( n14184 , n6770 );
    not g16076 ( n7986 , n30331 );
    xnor g16077 ( n16493 , n15717 , n151 );
    xnor g16078 ( n24524 , n4950 , n23218 );
    not g16079 ( n1829 , n7435 );
    and g16080 ( n30496 , n638 , n15611 );
    xnor g16081 ( n20841 , n25699 , n17051 );
    xor g16082 ( n25350 , n153 , n26848 );
    not g16083 ( n8292 , n22675 );
    and g16084 ( n11904 , n31322 , n19698 );
    nor g16085 ( n6466 , n30887 , n28983 );
    and g16086 ( n14783 , n26651 , n9541 );
    and g16087 ( n7260 , n10422 , n15775 );
    not g16088 ( n2174 , n17729 );
    not g16089 ( n1355 , n7173 );
    not g16090 ( n24918 , n7583 );
    not g16091 ( n12091 , n31655 );
    nor g16092 ( n12490 , n12429 , n14000 );
    nor g16093 ( n17571 , n13939 , n10938 );
    not g16094 ( n10757 , n17644 );
    or g16095 ( n5244 , n13269 , n4681 );
    xnor g16096 ( n21320 , n29826 , n5082 );
    not g16097 ( n26390 , n22660 );
    and g16098 ( n14729 , n16906 , n31387 );
    not g16099 ( n17085 , n853 );
    xnor g16100 ( n24770 , n10811 , n6550 );
    nor g16101 ( n2011 , n10376 , n12320 );
    not g16102 ( n14467 , n2477 );
    not g16103 ( n2319 , n28372 );
    or g16104 ( n501 , n4560 , n3118 );
    or g16105 ( n31172 , n30344 , n11184 );
    not g16106 ( n20403 , n26343 );
    or g16107 ( n7501 , n6984 , n30349 );
    or g16108 ( n2816 , n21607 , n23437 );
    or g16109 ( n27158 , n24437 , n10608 );
    xnor g16110 ( n20238 , n19185 , n11361 );
    not g16111 ( n23045 , n29279 );
    not g16112 ( n23657 , n6165 );
    xnor g16113 ( n30169 , n11655 , n209 );
    not g16114 ( n14827 , n21863 );
    or g16115 ( n1474 , n21640 , n25772 );
    xnor g16116 ( n27381 , n17410 , n16950 );
    not g16117 ( n3056 , n8185 );
    or g16118 ( n21512 , n15914 , n10515 );
    xnor g16119 ( n9797 , n22981 , n26193 );
    or g16120 ( n10170 , n31578 , n27125 );
    xnor g16121 ( n7694 , n26006 , n29249 );
    xnor g16122 ( n19207 , n25710 , n292 );
    xnor g16123 ( n6254 , n266 , n16938 );
    xnor g16124 ( n29057 , n15588 , n16075 );
    xnor g16125 ( n12805 , n30963 , n20084 );
    or g16126 ( n15304 , n13670 , n12414 );
    or g16127 ( n2361 , n14437 , n9730 );
    not g16128 ( n21208 , n6445 );
    and g16129 ( n31816 , n26113 , n19389 );
    not g16130 ( n17428 , n17599 );
    not g16131 ( n16719 , n12246 );
    and g16132 ( n10727 , n18520 , n12718 );
    xnor g16133 ( n22304 , n25355 , n21209 );
    xnor g16134 ( n8790 , n4192 , n15170 );
    not g16135 ( n30691 , n20905 );
    not g16136 ( n12910 , n740 );
    or g16137 ( n6675 , n1317 , n15629 );
    or g16138 ( n16074 , n8901 , n20883 );
    not g16139 ( n14961 , n6399 );
    not g16140 ( n25145 , n24710 );
    or g16141 ( n6312 , n17459 , n24863 );
    and g16142 ( n15282 , n11647 , n5557 );
    not g16143 ( n7160 , n14527 );
    nor g16144 ( n17949 , n28198 , n13597 );
    xnor g16145 ( n26355 , n2963 , n9239 );
    or g16146 ( n9672 , n21122 , n6253 );
    or g16147 ( n20247 , n16794 , n21687 );
    xor g16148 ( n690 , n15053 , n7520 );
    xnor g16149 ( n2788 , n14013 , n29844 );
    not g16150 ( n1463 , n6137 );
    and g16151 ( n9298 , n12005 , n11135 );
    nor g16152 ( n22910 , n26235 , n20187 );
    not g16153 ( n25827 , n12803 );
    not g16154 ( n19765 , n15519 );
    not g16155 ( n7876 , n20332 );
    not g16156 ( n27317 , n22292 );
    not g16157 ( n1270 , n9565 );
    not g16158 ( n22043 , n6449 );
    and g16159 ( n9899 , n663 , n18320 );
    xnor g16160 ( n8798 , n9097 , n17173 );
    or g16161 ( n1321 , n2782 , n27979 );
    not g16162 ( n3588 , n2231 );
    nor g16163 ( n26594 , n25871 , n18975 );
    not g16164 ( n25175 , n27357 );
    and g16165 ( n6051 , n9979 , n20401 );
    or g16166 ( n4816 , n369 , n26895 );
    or g16167 ( n14540 , n21327 , n1508 );
    xnor g16168 ( n21730 , n10221 , n3040 );
    and g16169 ( n17365 , n10945 , n2790 );
    not g16170 ( n17496 , n15010 );
    or g16171 ( n21775 , n11893 , n12848 );
    xnor g16172 ( n28750 , n12457 , n6591 );
    xnor g16173 ( n12017 , n30277 , n13599 );
    and g16174 ( n17694 , n5039 , n18099 );
    xnor g16175 ( n3895 , n13057 , n10210 );
    and g16176 ( n5946 , n16378 , n16107 );
    nor g16177 ( n14514 , n18028 , n4467 );
    or g16178 ( n15455 , n13776 , n9109 );
    xnor g16179 ( n8876 , n10660 , n23012 );
    not g16180 ( n23701 , n27238 );
    and g16181 ( n3945 , n11580 , n22845 );
    and g16182 ( n8216 , n12592 , n22735 );
    xnor g16183 ( n5908 , n8817 , n13681 );
    not g16184 ( n2808 , n18370 );
    not g16185 ( n13768 , n22325 );
    nor g16186 ( n7920 , n810 , n31076 );
    not g16187 ( n678 , n30180 );
    or g16188 ( n24887 , n8418 , n6046 );
    or g16189 ( n23631 , n2188 , n27785 );
    not g16190 ( n1979 , n12986 );
    or g16191 ( n13847 , n4658 , n29542 );
    or g16192 ( n14071 , n16406 , n8863 );
    or g16193 ( n22231 , n6957 , n28226 );
    or g16194 ( n5587 , n7146 , n29254 );
    and g16195 ( n3560 , n26124 , n15657 );
    xnor g16196 ( n25370 , n6172 , n22316 );
    and g16197 ( n26341 , n14879 , n15233 );
    xnor g16198 ( n18904 , n16122 , n16599 );
    or g16199 ( n20081 , n15468 , n27289 );
    not g16200 ( n6901 , n18155 );
    not g16201 ( n25374 , n7414 );
    xnor g16202 ( n12974 , n24313 , n28494 );
    or g16203 ( n11562 , n19958 , n22084 );
    not g16204 ( n21982 , n10909 );
    xnor g16205 ( n4193 , n29772 , n9590 );
    nor g16206 ( n15071 , n13473 , n13594 );
    xnor g16207 ( n1059 , n7052 , n16193 );
    or g16208 ( n972 , n28300 , n30501 );
    not g16209 ( n24353 , n26549 );
    or g16210 ( n17513 , n21838 , n18089 );
    or g16211 ( n16358 , n25760 , n28527 );
    xnor g16212 ( n1882 , n19905 , n8609 );
    not g16213 ( n1800 , n7626 );
    not g16214 ( n289 , n24132 );
    and g16215 ( n24009 , n8136 , n22063 );
    or g16216 ( n11240 , n23350 , n737 );
    not g16217 ( n6962 , n23632 );
    not g16218 ( n11667 , n4759 );
    xnor g16219 ( n4647 , n4101 , n12858 );
    xnor g16220 ( n379 , n20349 , n24081 );
    or g16221 ( n432 , n18219 , n5549 );
    not g16222 ( n18503 , n30458 );
    and g16223 ( n9676 , n13699 , n20248 );
    or g16224 ( n17442 , n21312 , n24989 );
    nor g16225 ( n13305 , n22451 , n10504 );
    and g16226 ( n24550 , n9903 , n6420 );
    xnor g16227 ( n28993 , n23480 , n21625 );
    and g16228 ( n21854 , n16863 , n13470 );
    xnor g16229 ( n27031 , n17114 , n10447 );
    and g16230 ( n940 , n6410 , n28339 );
    not g16231 ( n20289 , n3810 );
    xnor g16232 ( n20587 , n16967 , n1494 );
    xnor g16233 ( n25603 , n10240 , n9762 );
    nor g16234 ( n9515 , n26904 , n19437 );
    nor g16235 ( n14684 , n31204 , n4744 );
    or g16236 ( n31833 , n30980 , n7454 );
    and g16237 ( n16048 , n5738 , n28153 );
    not g16238 ( n17841 , n1293 );
    and g16239 ( n10762 , n5480 , n12426 );
    and g16240 ( n7365 , n14104 , n31896 );
    xnor g16241 ( n14008 , n19387 , n6407 );
    not g16242 ( n7646 , n15447 );
    not g16243 ( n31211 , n18940 );
    not g16244 ( n27816 , n25878 );
    nor g16245 ( n504 , n18652 , n27747 );
    not g16246 ( n2870 , n18983 );
    nor g16247 ( n19601 , n7180 , n493 );
    or g16248 ( n17203 , n4788 , n76 );
    not g16249 ( n31585 , n18723 );
    or g16250 ( n23517 , n4890 , n20505 );
    or g16251 ( n10875 , n29392 , n10183 );
    nor g16252 ( n7955 , n10888 , n24457 );
    or g16253 ( n2186 , n32003 , n23587 );
    not g16254 ( n11737 , n19315 );
    or g16255 ( n25892 , n529 , n5234 );
    xnor g16256 ( n30364 , n12011 , n24266 );
    and g16257 ( n5412 , n24385 , n20055 );
    not g16258 ( n2457 , n20315 );
    nor g16259 ( n17655 , n21136 , n31366 );
    not g16260 ( n25496 , n17960 );
    xnor g16261 ( n9352 , n20432 , n4027 );
    xnor g16262 ( n179 , n30668 , n12242 );
    not g16263 ( n18485 , n9342 );
    not g16264 ( n14450 , n28288 );
    xnor g16265 ( n1974 , n793 , n20815 );
    or g16266 ( n26384 , n18838 , n30500 );
    and g16267 ( n10330 , n1237 , n17309 );
    or g16268 ( n25992 , n21354 , n5597 );
    or g16269 ( n27945 , n891 , n22203 );
    and g16270 ( n14645 , n5910 , n2988 );
    xnor g16271 ( n15665 , n25793 , n24137 );
    or g16272 ( n21022 , n7793 , n6379 );
    or g16273 ( n4369 , n685 , n18407 );
    and g16274 ( n31458 , n28063 , n14802 );
    xnor g16275 ( n9883 , n17095 , n19405 );
    or g16276 ( n6220 , n11174 , n20188 );
    xnor g16277 ( n23771 , n4430 , n13615 );
    xnor g16278 ( n31396 , n18111 , n24829 );
    not g16279 ( n26689 , n19801 );
    not g16280 ( n3804 , n31878 );
    and g16281 ( n1240 , n27232 , n10054 );
    or g16282 ( n4878 , n16609 , n5402 );
    xnor g16283 ( n18372 , n1711 , n18367 );
    not g16284 ( n5391 , n29162 );
    not g16285 ( n25035 , n18124 );
    xnor g16286 ( n448 , n23033 , n6669 );
    or g16287 ( n28042 , n11228 , n15856 );
    xnor g16288 ( n22509 , n3787 , n12312 );
    nor g16289 ( n26737 , n6704 , n26846 );
    not g16290 ( n16459 , n15429 );
    or g16291 ( n5803 , n24034 , n23439 );
    not g16292 ( n1125 , n7675 );
    not g16293 ( n2537 , n28112 );
    not g16294 ( n18192 , n29567 );
    and g16295 ( n5420 , n21472 , n31600 );
    and g16296 ( n28839 , n5795 , n11179 );
    not g16297 ( n16958 , n30913 );
    not g16298 ( n6653 , n2542 );
    or g16299 ( n4980 , n15631 , n12482 );
    not g16300 ( n14386 , n25295 );
    xnor g16301 ( n7005 , n9116 , n7210 );
    not g16302 ( n27670 , n9825 );
    and g16303 ( n9178 , n31103 , n4442 );
    not g16304 ( n11785 , n17867 );
    xnor g16305 ( n20772 , n26712 , n30692 );
    xnor g16306 ( n16822 , n493 , n7180 );
    xnor g16307 ( n28615 , n21997 , n7068 );
    xnor g16308 ( n21237 , n1057 , n3108 );
    not g16309 ( n4065 , n8030 );
    not g16310 ( n14390 , n23047 );
    and g16311 ( n4455 , n24763 , n3188 );
    not g16312 ( n1530 , n5360 );
    and g16313 ( n8946 , n16589 , n224 );
    and g16314 ( n31909 , n24541 , n19148 );
    or g16315 ( n25544 , n26532 , n10502 );
    not g16316 ( n1212 , n29349 );
    not g16317 ( n18177 , n8848 );
    not g16318 ( n23817 , n30405 );
    nor g16319 ( n14330 , n21671 , n31479 );
    and g16320 ( n21226 , n13014 , n5321 );
    not g16321 ( n6756 , n4942 );
    or g16322 ( n4902 , n15227 , n11274 );
    and g16323 ( n29267 , n31061 , n10297 );
    not g16324 ( n17969 , n25173 );
    not g16325 ( n17382 , n24070 );
    xnor g16326 ( n22527 , n29766 , n11368 );
    and g16327 ( n30415 , n8156 , n15918 );
    not g16328 ( n17913 , n2064 );
    and g16329 ( n19096 , n6503 , n1553 );
    or g16330 ( n14151 , n4341 , n24183 );
    xnor g16331 ( n31144 , n8216 , n4177 );
    and g16332 ( n29481 , n24754 , n25433 );
    nor g16333 ( n1464 , n4878 , n883 );
    or g16334 ( n18174 , n27229 , n11854 );
    and g16335 ( n15867 , n16636 , n24119 );
    or g16336 ( n21517 , n8424 , n11858 );
    and g16337 ( n15317 , n23866 , n25535 );
    or g16338 ( n12868 , n14431 , n6485 );
    not g16339 ( n14346 , n16541 );
    or g16340 ( n19784 , n22933 , n16419 );
    or g16341 ( n14193 , n32014 , n28309 );
    not g16342 ( n20655 , n100 );
    and g16343 ( n7001 , n6380 , n31226 );
    nor g16344 ( n24587 , n9338 , n7379 );
    or g16345 ( n13126 , n23770 , n559 );
    buf g16346 ( n22294 , n14392 );
    or g16347 ( n9074 , n21829 , n9280 );
    not g16348 ( n12781 , n4120 );
    and g16349 ( n1510 , n1110 , n25645 );
    xnor g16350 ( n15416 , n16224 , n15783 );
    or g16351 ( n7782 , n131 , n28077 );
    or g16352 ( n27987 , n1077 , n26299 );
    or g16353 ( n21860 , n25739 , n3237 );
    and g16354 ( n13904 , n21913 , n14529 );
    xnor g16355 ( n12943 , n705 , n2175 );
    or g16356 ( n25134 , n7226 , n14261 );
    not g16357 ( n17893 , n6322 );
    xnor g16358 ( n22270 , n21732 , n3547 );
    xnor g16359 ( n26178 , n17223 , n8298 );
    not g16360 ( n20046 , n20864 );
    and g16361 ( n16188 , n2769 , n27281 );
    xnor g16362 ( n14907 , n11073 , n31042 );
    not g16363 ( n21934 , n8944 );
    xnor g16364 ( n28474 , n10589 , n16660 );
    or g16365 ( n17951 , n6609 , n13923 );
    or g16366 ( n5199 , n30495 , n10900 );
    not g16367 ( n13698 , n19557 );
    not g16368 ( n20187 , n3080 );
    not g16369 ( n5406 , n2562 );
    xnor g16370 ( n25978 , n25116 , n19038 );
    or g16371 ( n11336 , n10737 , n30419 );
    nor g16372 ( n10412 , n24785 , n5535 );
    not g16373 ( n26586 , n21572 );
    or g16374 ( n4634 , n4627 , n19997 );
    xnor g16375 ( n29741 , n23234 , n2381 );
    xnor g16376 ( n25630 , n5908 , n20359 );
    or g16377 ( n2493 , n31152 , n6827 );
    nor g16378 ( n8809 , n9939 , n9524 );
    xnor g16379 ( n5499 , n30002 , n9655 );
    and g16380 ( n27515 , n31180 , n29549 );
    xor g16381 ( n11059 , n30356 , n19393 );
    xnor g16382 ( n22013 , n14711 , n6534 );
    and g16383 ( n9243 , n11560 , n26390 );
    xnor g16384 ( n20394 , n4240 , n31722 );
    xnor g16385 ( n14148 , n17459 , n13184 );
    and g16386 ( n2969 , n13886 , n13043 );
    nor g16387 ( n19985 , n11648 , n19979 );
    nor g16388 ( n8541 , n2688 , n12610 );
    not g16389 ( n21263 , n6492 );
    not g16390 ( n21528 , n22844 );
    xnor g16391 ( n29545 , n29427 , n2337 );
    or g16392 ( n20617 , n11749 , n12058 );
    xnor g16393 ( n6976 , n10480 , n29006 );
    not g16394 ( n8080 , n3532 );
    xnor g16395 ( n9800 , n19854 , n21170 );
    and g16396 ( n18427 , n28913 , n8919 );
    xnor g16397 ( n11982 , n11223 , n20175 );
    and g16398 ( n16823 , n1904 , n9848 );
    or g16399 ( n500 , n1095 , n8451 );
    not g16400 ( n15198 , n2058 );
    not g16401 ( n15852 , n20861 );
    not g16402 ( n110 , n13434 );
    or g16403 ( n27884 , n29158 , n24869 );
    and g16404 ( n28172 , n25595 , n18534 );
    nor g16405 ( n3441 , n18002 , n4618 );
    or g16406 ( n3126 , n18054 , n26098 );
    or g16407 ( n2593 , n13129 , n27216 );
    xnor g16408 ( n19534 , n15528 , n19518 );
    not g16409 ( n4157 , n27454 );
    and g16410 ( n10760 , n12919 , n32027 );
    or g16411 ( n2988 , n7757 , n15648 );
    not g16412 ( n7504 , n29109 );
    xnor g16413 ( n13596 , n17799 , n11969 );
    xnor g16414 ( n20011 , n24447 , n20022 );
    nor g16415 ( n17244 , n16312 , n3473 );
    xor g16416 ( n24614 , n9498 , n14670 );
    xnor g16417 ( n29951 , n21438 , n8632 );
    not g16418 ( n20490 , n12756 );
    not g16419 ( n4964 , n11271 );
    xnor g16420 ( n4661 , n6166 , n12971 );
    xnor g16421 ( n15186 , n30183 , n23663 );
    and g16422 ( n21097 , n21527 , n6791 );
    not g16423 ( n20943 , n15151 );
    and g16424 ( n31158 , n25725 , n16496 );
    or g16425 ( n15695 , n17457 , n3661 );
    not g16426 ( n25532 , n7787 );
    not g16427 ( n19252 , n15923 );
    not g16428 ( n9726 , n21425 );
    and g16429 ( n14509 , n7227 , n11352 );
    and g16430 ( n30878 , n5263 , n16332 );
    not g16431 ( n30998 , n18572 );
    nor g16432 ( n6989 , n7355 , n13949 );
    xnor g16433 ( n8168 , n12802 , n775 );
    xnor g16434 ( n1571 , n28052 , n16869 );
    or g16435 ( n31706 , n2274 , n5590 );
    and g16436 ( n19872 , n19329 , n1834 );
    or g16437 ( n5776 , n914 , n920 );
    and g16438 ( n26712 , n20265 , n3018 );
    nor g16439 ( n10991 , n11361 , n10837 );
    xnor g16440 ( n21809 , n31448 , n11984 );
    not g16441 ( n14785 , n19161 );
    nor g16442 ( n2110 , n13978 , n28264 );
    not g16443 ( n12319 , n5747 );
    or g16444 ( n15250 , n17027 , n22897 );
    xnor g16445 ( n22733 , n21261 , n3076 );
    not g16446 ( n19384 , n6808 );
    xnor g16447 ( n29171 , n123 , n25065 );
    not g16448 ( n23059 , n16987 );
    not g16449 ( n25445 , n2998 );
    or g16450 ( n3493 , n21381 , n26931 );
    not g16451 ( n12882 , n6331 );
    not g16452 ( n21565 , n25067 );
    not g16453 ( n3491 , n30105 );
    not g16454 ( n30255 , n25837 );
    or g16455 ( n2158 , n6581 , n2203 );
    or g16456 ( n25949 , n15346 , n22885 );
    not g16457 ( n14688 , n3516 );
    not g16458 ( n10814 , n12683 );
    not g16459 ( n1512 , n9209 );
    not g16460 ( n31388 , n6666 );
    or g16461 ( n29608 , n23620 , n31813 );
    xnor g16462 ( n30889 , n3765 , n2963 );
    not g16463 ( n23826 , n20905 );
    or g16464 ( n4559 , n10887 , n17443 );
    xnor g16465 ( n23360 , n17662 , n4891 );
    and g16466 ( n4724 , n30125 , n13637 );
    xnor g16467 ( n4810 , n7375 , n20098 );
    not g16468 ( n4542 , n25871 );
    nor g16469 ( n10340 , n5069 , n28857 );
    or g16470 ( n27392 , n17332 , n19089 );
    xnor g16471 ( n14677 , n1048 , n5388 );
    and g16472 ( n6343 , n23430 , n19524 );
    xnor g16473 ( n12861 , n24465 , n30956 );
    not g16474 ( n6528 , n14427 );
    or g16475 ( n22196 , n20991 , n12456 );
    nor g16476 ( n30683 , n27440 , n5425 );
    not g16477 ( n12305 , n20050 );
    nor g16478 ( n978 , n9657 , n5399 );
    and g16479 ( n22272 , n25921 , n9672 );
    not g16480 ( n900 , n17622 );
    nor g16481 ( n26879 , n22746 , n20420 );
    or g16482 ( n13115 , n7500 , n22463 );
    nor g16483 ( n31555 , n238 , n30565 );
    and g16484 ( n426 , n14360 , n8458 );
    not g16485 ( n31584 , n20726 );
    and g16486 ( n17443 , n2077 , n3054 );
    not g16487 ( n8348 , n30593 );
    not g16488 ( n26250 , n6691 );
    xnor g16489 ( n26362 , n24825 , n29980 );
    or g16490 ( n20099 , n26622 , n16380 );
    not g16491 ( n2718 , n29486 );
    xnor g16492 ( n20857 , n5549 , n7019 );
    or g16493 ( n26556 , n4253 , n1537 );
    and g16494 ( n5399 , n4565 , n1926 );
    xnor g16495 ( n30608 , n1891 , n27151 );
    not g16496 ( n18956 , n26424 );
    not g16497 ( n12131 , n10056 );
    xnor g16498 ( n12645 , n702 , n30940 );
    or g16499 ( n25131 , n15545 , n19383 );
    xnor g16500 ( n106 , n5149 , n16609 );
    and g16501 ( n14508 , n30752 , n19006 );
    xnor g16502 ( n27104 , n21124 , n15156 );
    xor g16503 ( n31193 , n21057 , n1339 );
    nor g16504 ( n2546 , n10799 , n687 );
    and g16505 ( n8229 , n5609 , n10136 );
    or g16506 ( n7176 , n2934 , n24773 );
    xnor g16507 ( n731 , n26962 , n9494 );
    xnor g16508 ( n19525 , n19585 , n30278 );
    or g16509 ( n23661 , n7186 , n3413 );
    xnor g16510 ( n16694 , n10540 , n3172 );
    xnor g16511 ( n4114 , n18645 , n23306 );
    xnor g16512 ( n2878 , n9346 , n6100 );
    xnor g16513 ( n19619 , n30507 , n3079 );
    xnor g16514 ( n20433 , n31826 , n2547 );
    not g16515 ( n30252 , n27774 );
    not g16516 ( n29224 , n28896 );
    or g16517 ( n22520 , n5530 , n9210 );
    and g16518 ( n17252 , n6519 , n6623 );
    or g16519 ( n19819 , n16998 , n17641 );
    xnor g16520 ( n7398 , n30792 , n10017 );
    or g16521 ( n19640 , n27431 , n2073 );
    not g16522 ( n2802 , n11651 );
    xnor g16523 ( n3145 , n13316 , n26080 );
    or g16524 ( n11508 , n8074 , n5191 );
    xnor g16525 ( n24748 , n3810 , n4847 );
    and g16526 ( n15497 , n13200 , n30130 );
    not g16527 ( n5573 , n28621 );
    xnor g16528 ( n8153 , n29801 , n26109 );
    xnor g16529 ( n10438 , n7815 , n10115 );
    xnor g16530 ( n23280 , n14147 , n11462 );
    not g16531 ( n9468 , n10386 );
    not g16532 ( n18127 , n9387 );
    or g16533 ( n11001 , n24020 , n17377 );
    not g16534 ( n10493 , n11288 );
    or g16535 ( n10457 , n4278 , n21314 );
    or g16536 ( n26846 , n9600 , n8727 );
    xnor g16537 ( n19459 , n25610 , n2832 );
    and g16538 ( n18313 , n30050 , n29608 );
    not g16539 ( n29472 , n31204 );
    or g16540 ( n710 , n29941 , n3151 );
    xnor g16541 ( n6719 , n12114 , n16190 );
    not g16542 ( n25023 , n11519 );
    not g16543 ( n8394 , n17609 );
    or g16544 ( n4932 , n19313 , n15554 );
    xnor g16545 ( n16943 , n24854 , n4849 );
    xnor g16546 ( n396 , n27308 , n9352 );
    or g16547 ( n4407 , n15966 , n20682 );
    or g16548 ( n21907 , n6716 , n23880 );
    not g16549 ( n26992 , n22626 );
    not g16550 ( n22472 , n17661 );
    not g16551 ( n21663 , n3792 );
    xnor g16552 ( n27071 , n3322 , n3345 );
    not g16553 ( n17826 , n29949 );
    and g16554 ( n13095 , n15743 , n24684 );
    nor g16555 ( n19567 , n28555 , n12832 );
    or g16556 ( n14698 , n20055 , n20556 );
    or g16557 ( n30243 , n13464 , n2352 );
    and g16558 ( n11396 , n1654 , n28239 );
    and g16559 ( n31125 , n15861 , n21941 );
    not g16560 ( n16241 , n6026 );
    not g16561 ( n26148 , n8281 );
    xnor g16562 ( n10647 , n24683 , n4573 );
    xnor g16563 ( n25759 , n5989 , n15797 );
    or g16564 ( n24790 , n19181 , n11909 );
    xnor g16565 ( n14287 , n20340 , n29502 );
    and g16566 ( n29914 , n30782 , n32026 );
    and g16567 ( n26313 , n11100 , n4325 );
    and g16568 ( n9928 , n13060 , n11737 );
    and g16569 ( n28594 , n7099 , n4799 );
    xnor g16570 ( n17953 , n22888 , n30236 );
    xnor g16571 ( n30079 , n4113 , n27661 );
    or g16572 ( n14586 , n31567 , n4940 );
    xnor g16573 ( n28318 , n10139 , n25760 );
    and g16574 ( n17393 , n9272 , n941 );
    and g16575 ( n2063 , n16770 , n6918 );
    xnor g16576 ( n31711 , n27378 , n13074 );
    and g16577 ( n12636 , n1254 , n5813 );
    not g16578 ( n16744 , n22245 );
    or g16579 ( n18813 , n29480 , n8247 );
    and g16580 ( n354 , n11350 , n11846 );
    not g16581 ( n9195 , n26368 );
    and g16582 ( n23155 , n21650 , n13525 );
    not g16583 ( n23998 , n28165 );
    nor g16584 ( n31290 , n31301 , n6302 );
    xnor g16585 ( n3313 , n9094 , n28835 );
    and g16586 ( n21434 , n19994 , n26621 );
    and g16587 ( n26970 , n6635 , n18414 );
    not g16588 ( n30207 , n10158 );
    or g16589 ( n15728 , n3879 , n11366 );
    or g16590 ( n14921 , n22968 , n21137 );
    and g16591 ( n30077 , n17228 , n18183 );
    not g16592 ( n10542 , n22938 );
    or g16593 ( n31607 , n13416 , n16513 );
    not g16594 ( n17793 , n50 );
    or g16595 ( n29190 , n18841 , n22837 );
    xor g16596 ( n8764 , n12372 , n20135 );
    and g16597 ( n29561 , n16144 , n10450 );
    or g16598 ( n640 , n9095 , n16472 );
    or g16599 ( n9278 , n26351 , n19510 );
    xnor g16600 ( n21474 , n19132 , n508 );
    and g16601 ( n22789 , n12420 , n7176 );
    not g16602 ( n3025 , n20714 );
    xnor g16603 ( n19 , n1720 , n13635 );
    or g16604 ( n8899 , n19616 , n9397 );
    xnor g16605 ( n19268 , n14951 , n756 );
    or g16606 ( n6385 , n21110 , n498 );
    or g16607 ( n29425 , n14663 , n24313 );
    xnor g16608 ( n27988 , n10139 , n107 );
    not g16609 ( n5586 , n899 );
    and g16610 ( n25088 , n7935 , n31161 );
    not g16611 ( n3332 , n28742 );
    and g16612 ( n14829 , n21347 , n14486 );
    xnor g16613 ( n23104 , n1195 , n15178 );
    not g16614 ( n2648 , n5494 );
    or g16615 ( n16220 , n18363 , n15923 );
    not g16616 ( n8781 , n28878 );
    xnor g16617 ( n17875 , n10139 , n238 );
    and g16618 ( n25795 , n16063 , n10184 );
    and g16619 ( n21946 , n6897 , n8614 );
    not g16620 ( n8421 , n31323 );
    not g16621 ( n2516 , n14317 );
    not g16622 ( n1859 , n7661 );
    and g16623 ( n24942 , n17002 , n8336 );
    not g16624 ( n26122 , n19372 );
    and g16625 ( n14647 , n28784 , n18365 );
    xnor g16626 ( n14336 , n21189 , n15870 );
    or g16627 ( n4578 , n12905 , n21662 );
    and g16628 ( n27735 , n11141 , n24906 );
    xnor g16629 ( n13211 , n20140 , n15960 );
    not g16630 ( n20306 , n6714 );
    and g16631 ( n13574 , n26917 , n4923 );
    or g16632 ( n410 , n25274 , n23222 );
    xnor g16633 ( n9458 , n30024 , n9134 );
    or g16634 ( n21183 , n8620 , n24639 );
    xnor g16635 ( n9906 , n8550 , n29683 );
    or g16636 ( n15775 , n17116 , n7132 );
    and g16637 ( n14944 , n18798 , n22449 );
    not g16638 ( n11493 , n24214 );
    and g16639 ( n20936 , n11027 , n108 );
    or g16640 ( n17463 , n2234 , n18935 );
    not g16641 ( n23627 , n25391 );
    nor g16642 ( n20637 , n13957 , n24510 );
    xnor g16643 ( n1918 , n15865 , n20260 );
    or g16644 ( n27202 , n15402 , n8398 );
    buf g16645 ( n11851 , n24463 );
    not g16646 ( n3122 , n8317 );
    or g16647 ( n13623 , n17541 , n662 );
    not g16648 ( n16523 , n5374 );
    xnor g16649 ( n29317 , n8640 , n32020 );
    or g16650 ( n4331 , n19624 , n14539 );
    xnor g16651 ( n16140 , n31497 , n23380 );
    or g16652 ( n16990 , n12173 , n25484 );
    xnor g16653 ( n29266 , n1077 , n19283 );
    not g16654 ( n2767 , n26182 );
    nor g16655 ( n31559 , n25997 , n20408 );
    xor g16656 ( n6136 , n16208 , n23727 );
    nor g16657 ( n6038 , n30228 , n15485 );
    not g16658 ( n22047 , n31960 );
    not g16659 ( n17688 , n1725 );
    or g16660 ( n5282 , n2112 , n16331 );
    not g16661 ( n26724 , n31655 );
    xnor g16662 ( n12960 , n3553 , n899 );
    and g16663 ( n24877 , n215 , n12364 );
    or g16664 ( n181 , n11643 , n8802 );
    xnor g16665 ( n5706 , n19653 , n26355 );
    not g16666 ( n26184 , n18989 );
    not g16667 ( n16720 , n12493 );
    or g16668 ( n31699 , n16498 , n16520 );
    xnor g16669 ( n20105 , n9476 , n14112 );
    not g16670 ( n447 , n27851 );
    not g16671 ( n6416 , n20038 );
    nor g16672 ( n16567 , n10109 , n13704 );
    not g16673 ( n30277 , n16068 );
    or g16674 ( n5308 , n17986 , n13548 );
    not g16675 ( n129 , n22814 );
    xnor g16676 ( n24937 , n103 , n10823 );
    not g16677 ( n19023 , n14962 );
    xnor g16678 ( n18211 , n4025 , n24938 );
    not g16679 ( n274 , n31038 );
    not g16680 ( n16638 , n9803 );
    not g16681 ( n3725 , n23145 );
    xnor g16682 ( n13813 , n6214 , n12455 );
    not g16683 ( n22688 , n831 );
    or g16684 ( n5669 , n295 , n29035 );
    nor g16685 ( n27279 , n3810 , n25794 );
    or g16686 ( n31025 , n31187 , n22966 );
    xnor g16687 ( n11611 , n23067 , n1935 );
    and g16688 ( n26845 , n16 , n7927 );
    nor g16689 ( n19429 , n13145 , n12198 );
    nor g16690 ( n18677 , n22867 , n2734 );
    xor g16691 ( n20916 , n9337 , n29293 );
    not g16692 ( n24247 , n19432 );
    or g16693 ( n6692 , n9185 , n19892 );
    not g16694 ( n28907 , n2323 );
    nor g16695 ( n1005 , n17417 , n20289 );
    or g16696 ( n11875 , n3750 , n5970 );
    and g16697 ( n9738 , n1156 , n25473 );
    and g16698 ( n23845 , n2897 , n28118 );
    not g16699 ( n25106 , n23046 );
    xnor g16700 ( n29 , n21590 , n6183 );
    or g16701 ( n28228 , n23603 , n3124 );
    xnor g16702 ( n22120 , n12770 , n9967 );
    not g16703 ( n8800 , n17127 );
    and g16704 ( n595 , n5648 , n15086 );
    and g16705 ( n9503 , n7092 , n19003 );
    not g16706 ( n20441 , n14949 );
    or g16707 ( n27620 , n19913 , n28674 );
    and g16708 ( n16219 , n17020 , n15974 );
    xnor g16709 ( n13780 , n6428 , n31111 );
    and g16710 ( n7805 , n13168 , n27989 );
    xnor g16711 ( n24449 , n27619 , n19237 );
    buf g16712 ( n11581 , n21923 );
    not g16713 ( n11861 , n30971 );
    not g16714 ( n6247 , n28818 );
    xnor g16715 ( n16290 , n23195 , n13700 );
    not g16716 ( n31511 , n15254 );
    or g16717 ( n21200 , n11132 , n24344 );
    not g16718 ( n30901 , n26100 );
    or g16719 ( n5761 , n24903 , n28840 );
    and g16720 ( n326 , n28306 , n31918 );
    or g16721 ( n23386 , n12403 , n15450 );
    and g16722 ( n15957 , n28336 , n31203 );
    xnor g16723 ( n1292 , n24599 , n29292 );
    and g16724 ( n11499 , n5699 , n11785 );
    and g16725 ( n28186 , n27526 , n16074 );
    nor g16726 ( n11713 , n20108 , n22574 );
    nor g16727 ( n31018 , n12777 , n31851 );
    xnor g16728 ( n16250 , n20100 , n30605 );
    not g16729 ( n24890 , n32020 );
    or g16730 ( n19565 , n26359 , n12439 );
    not g16731 ( n7380 , n11816 );
    nor g16732 ( n7399 , n20210 , n25758 );
    xnor g16733 ( n764 , n12459 , n23255 );
    or g16734 ( n24915 , n9064 , n10366 );
    not g16735 ( n588 , n13220 );
    or g16736 ( n24146 , n22173 , n29844 );
    xnor g16737 ( n8245 , n6481 , n3312 );
    and g16738 ( n21054 , n8871 , n9804 );
    not g16739 ( n8220 , n10947 );
    or g16740 ( n2750 , n28853 , n12047 );
    xnor g16741 ( n13141 , n24905 , n18582 );
    and g16742 ( n19086 , n24367 , n8115 );
    xnor g16743 ( n2095 , n20188 , n13028 );
    xnor g16744 ( n24345 , n614 , n31481 );
    not g16745 ( n26988 , n26598 );
    or g16746 ( n24693 , n18578 , n15480 );
    nor g16747 ( n31381 , n8512 , n19768 );
    not g16748 ( n29945 , n31343 );
    or g16749 ( n31220 , n31649 , n14412 );
    not g16750 ( n4030 , n30703 );
    and g16751 ( n11819 , n3868 , n18603 );
    not g16752 ( n11440 , n16725 );
    xnor g16753 ( n7083 , n22765 , n23960 );
    xnor g16754 ( n32024 , n28308 , n8856 );
    not g16755 ( n15195 , n25421 );
    not g16756 ( n16208 , n2883 );
    not g16757 ( n17686 , n19328 );
    and g16758 ( n31732 , n1316 , n22533 );
    xnor g16759 ( n18135 , n3389 , n19255 );
    or g16760 ( n29485 , n11452 , n16307 );
    nor g16761 ( n9855 , n12998 , n1349 );
    nor g16762 ( n29022 , n6957 , n23088 );
    nor g16763 ( n14697 , n22550 , n7313 );
    not g16764 ( n6072 , n29615 );
    or g16765 ( n4901 , n1099 , n21414 );
    not g16766 ( n8641 , n8083 );
    not g16767 ( n21055 , n7434 );
    or g16768 ( n15754 , n7655 , n14604 );
    not g16769 ( n28824 , n19538 );
    and g16770 ( n21587 , n18162 , n11129 );
    xor g16771 ( n863 , n8348 , n27122 );
    or g16772 ( n30952 , n23195 , n10433 );
    nor g16773 ( n13290 , n1474 , n1727 );
    xnor g16774 ( n30239 , n12429 , n11305 );
    and g16775 ( n10216 , n18820 , n20881 );
    xor g16776 ( n10028 , n23710 , n29790 );
    xnor g16777 ( n10319 , n23999 , n17243 );
    or g16778 ( n31463 , n29283 , n27755 );
    or g16779 ( n28290 , n21485 , n29053 );
    or g16780 ( n13324 , n21774 , n10839 );
    not g16781 ( n8989 , n4057 );
    nor g16782 ( n5911 , n31411 , n9895 );
    or g16783 ( n9127 , n26020 , n22215 );
    xnor g16784 ( n11062 , n5491 , n28067 );
    not g16785 ( n2510 , n20198 );
    not g16786 ( n26590 , n17038 );
    and g16787 ( n29280 , n17671 , n10459 );
    or g16788 ( n19365 , n84 , n14241 );
    not g16789 ( n5869 , n20310 );
    or g16790 ( n14559 , n27881 , n21594 );
    xnor g16791 ( n11185 , n10214 , n27381 );
    nor g16792 ( n19831 , n17046 , n15940 );
    not g16793 ( n9784 , n3903 );
    nor g16794 ( n30408 , n17036 , n3967 );
    xnor g16795 ( n18052 , n7360 , n4090 );
    buf g16796 ( n10847 , n13971 );
    or g16797 ( n28954 , n17320 , n13905 );
    not g16798 ( n7659 , n21425 );
    nor g16799 ( n26096 , n30158 , n10514 );
    or g16800 ( n3024 , n25408 , n569 );
    and g16801 ( n2073 , n29268 , n28726 );
    not g16802 ( n18549 , n5071 );
    or g16803 ( n5807 , n1988 , n7829 );
    nor g16804 ( n25849 , n10034 , n17142 );
    not g16805 ( n14260 , n13092 );
    nor g16806 ( n1847 , n26996 , n11065 );
    and g16807 ( n2209 , n25702 , n16370 );
    not g16808 ( n1841 , n14872 );
    not g16809 ( n24615 , n11712 );
    or g16810 ( n5424 , n11297 , n8499 );
    xnor g16811 ( n18678 , n27163 , n6071 );
    xnor g16812 ( n25897 , n16547 , n1242 );
    not g16813 ( n18737 , n15064 );
    nor g16814 ( n3360 , n11143 , n13658 );
    nor g16815 ( n13097 , n8996 , n19506 );
    xnor g16816 ( n9898 , n5437 , n17316 );
    not g16817 ( n28322 , n320 );
    or g16818 ( n29644 , n21484 , n13443 );
    or g16819 ( n11739 , n23611 , n14332 );
    nor g16820 ( n24301 , n10928 , n900 );
    not g16821 ( n20760 , n31060 );
    not g16822 ( n848 , n4086 );
    or g16823 ( n3031 , n7593 , n25137 );
    xnor g16824 ( n28675 , n2704 , n8260 );
    xnor g16825 ( n26526 , n20421 , n31836 );
    nor g16826 ( n7340 , n10356 , n22232 );
    not g16827 ( n18070 , n29897 );
    nor g16828 ( n21357 , n28158 , n3759 );
    not g16829 ( n1654 , n28518 );
    not g16830 ( n14403 , n2469 );
    xnor g16831 ( n1226 , n9440 , n20966 );
    or g16832 ( n17167 , n13488 , n17536 );
    xnor g16833 ( n28752 , n28410 , n990 );
    and g16834 ( n28665 , n14662 , n17436 );
    and g16835 ( n24967 , n11066 , n18176 );
    xnor g16836 ( n11265 , n27137 , n11873 );
    not g16837 ( n11913 , n27670 );
    or g16838 ( n21123 , n28983 , n29397 );
    xnor g16839 ( n3764 , n10260 , n8051 );
    xnor g16840 ( n5458 , n10137 , n30739 );
    or g16841 ( n8663 , n12214 , n5306 );
    or g16842 ( n25706 , n23594 , n29147 );
    and g16843 ( n9094 , n28708 , n26538 );
    and g16844 ( n23063 , n26627 , n26758 );
    or g16845 ( n8709 , n27025 , n8412 );
    xnor g16846 ( n13654 , n27415 , n7343 );
    not g16847 ( n23074 , n17902 );
    and g16848 ( n30500 , n7963 , n31157 );
    xnor g16849 ( n19476 , n15777 , n23389 );
    or g16850 ( n29677 , n20128 , n26662 );
    nor g16851 ( n14908 , n24120 , n5270 );
    xnor g16852 ( n24530 , n12035 , n7314 );
    not g16853 ( n24068 , n12920 );
    and g16854 ( n24092 , n12219 , n7666 );
    not g16855 ( n19832 , n20317 );
    xnor g16856 ( n8082 , n31551 , n21142 );
    and g16857 ( n13776 , n794 , n12627 );
    and g16858 ( n16580 , n2905 , n27383 );
    or g16859 ( n20131 , n7354 , n29087 );
    or g16860 ( n24886 , n18558 , n10501 );
    not g16861 ( n26610 , n1236 );
    and g16862 ( n5790 , n23139 , n18787 );
    or g16863 ( n11602 , n31577 , n18323 );
    not g16864 ( n15111 , n14993 );
    nor g16865 ( n21364 , n19572 , n901 );
    or g16866 ( n22869 , n8486 , n8968 );
    xnor g16867 ( n8824 , n27659 , n29054 );
    or g16868 ( n12846 , n29802 , n24933 );
    or g16869 ( n18540 , n31949 , n13304 );
    xnor g16870 ( n23551 , n896 , n8378 );
    or g16871 ( n3448 , n7401 , n12709 );
    or g16872 ( n20707 , n27635 , n18030 );
    or g16873 ( n24264 , n17241 , n4785 );
    xnor g16874 ( n810 , n17222 , n1773 );
    xnor g16875 ( n21032 , n21734 , n23025 );
    or g16876 ( n15295 , n29774 , n6750 );
    not g16877 ( n9359 , n21492 );
    not g16878 ( n24595 , n12816 );
    and g16879 ( n10387 , n12394 , n7056 );
    not g16880 ( n28929 , n4143 );
    xnor g16881 ( n19546 , n2874 , n14209 );
    and g16882 ( n1052 , n23332 , n21999 );
    xnor g16883 ( n459 , n24438 , n14996 );
    not g16884 ( n11026 , n8246 );
    not g16885 ( n4966 , n31688 );
    or g16886 ( n8568 , n18916 , n16715 );
    or g16887 ( n29394 , n5032 , n31477 );
    and g16888 ( n9086 , n2917 , n14522 );
    xnor g16889 ( n13545 , n7245 , n19106 );
    and g16890 ( n593 , n24635 , n14127 );
    xnor g16891 ( n26054 , n20578 , n26630 );
    or g16892 ( n6037 , n23643 , n11412 );
    or g16893 ( n31922 , n4491 , n13889 );
    not g16894 ( n21817 , n11308 );
    or g16895 ( n19145 , n1737 , n26667 );
    and g16896 ( n30202 , n3865 , n20004 );
    nor g16897 ( n12503 , n24118 , n8647 );
    and g16898 ( n29005 , n3059 , n24660 );
    or g16899 ( n27190 , n27780 , n15202 );
    not g16900 ( n12659 , n31232 );
    nor g16901 ( n9866 , n28634 , n29095 );
    xor g16902 ( n13618 , n29364 , n18348 );
    not g16903 ( n4067 , n27453 );
    nor g16904 ( n4399 , n1057 , n3108 );
    xnor g16905 ( n28340 , n10518 , n18658 );
    and g16906 ( n2415 , n28526 , n16490 );
    or g16907 ( n766 , n11847 , n23470 );
    xor g16908 ( n19062 , n17590 , n8097 );
    xnor g16909 ( n358 , n4730 , n21784 );
    nor g16910 ( n6581 , n15390 , n22743 );
    xnor g16911 ( n5760 , n29181 , n28367 );
    xnor g16912 ( n7479 , n26659 , n31591 );
    or g16913 ( n30824 , n25123 , n15194 );
    xnor g16914 ( n17444 , n336 , n21659 );
    not g16915 ( n20305 , n29705 );
    or g16916 ( n3132 , n18996 , n12883 );
    and g16917 ( n9457 , n4713 , n30406 );
    or g16918 ( n5266 , n11771 , n26316 );
    or g16919 ( n29554 , n16347 , n16847 );
    not g16920 ( n3436 , n14467 );
    xnor g16921 ( n9274 , n4332 , n6853 );
    and g16922 ( n5731 , n15656 , n3647 );
    not g16923 ( n2271 , n12652 );
    xor g16924 ( n16312 , n370 , n17033 );
    or g16925 ( n400 , n20261 , n23413 );
    or g16926 ( n8913 , n28025 , n23261 );
    xnor g16927 ( n31993 , n31314 , n18701 );
    and g16928 ( n29321 , n18760 , n14026 );
    xnor g16929 ( n16741 , n3052 , n2224 );
    xnor g16930 ( n1314 , n14395 , n11273 );
    not g16931 ( n11222 , n17641 );
    xnor g16932 ( n12404 , n18335 , n19707 );
    and g16933 ( n19893 , n17307 , n31938 );
    or g16934 ( n15123 , n26805 , n13869 );
    or g16935 ( n9012 , n23859 , n12225 );
    and g16936 ( n6797 , n20441 , n28619 );
    not g16937 ( n13260 , n20115 );
    xnor g16938 ( n3094 , n12998 , n13410 );
    not g16939 ( n20012 , n26735 );
    not g16940 ( n10502 , n3459 );
    or g16941 ( n31810 , n10914 , n22343 );
    or g16942 ( n11190 , n30902 , n22101 );
    or g16943 ( n19204 , n12557 , n18301 );
    or g16944 ( n3594 , n18394 , n21038 );
    and g16945 ( n11569 , n7477 , n24330 );
    not g16946 ( n4992 , n17835 );
    and g16947 ( n16001 , n22431 , n23395 );
    and g16948 ( n16809 , n13117 , n9065 );
    xor g16949 ( n9275 , n15254 , n9822 );
    not g16950 ( n23130 , n9690 );
    not g16951 ( n21178 , n13437 );
    not g16952 ( n5137 , n9412 );
    or g16953 ( n10080 , n28305 , n26433 );
    or g16954 ( n3669 , n4617 , n22592 );
    or g16955 ( n12921 , n12553 , n29012 );
    xnor g16956 ( n7411 , n12302 , n29076 );
    nor g16957 ( n14191 , n4113 , n29683 );
    or g16958 ( n31116 , n11886 , n28073 );
    not g16959 ( n31626 , n24354 );
    and g16960 ( n19684 , n23120 , n6688 );
    and g16961 ( n14002 , n12066 , n3782 );
    xnor g16962 ( n16401 , n11043 , n29252 );
    not g16963 ( n22382 , n17995 );
    xnor g16964 ( n3930 , n911 , n1115 );
    or g16965 ( n26132 , n2939 , n1590 );
    and g16966 ( n28353 , n6656 , n15313 );
    and g16967 ( n26699 , n16736 , n8264 );
    or g16968 ( n6677 , n16803 , n23342 );
    or g16969 ( n27057 , n13025 , n31158 );
    and g16970 ( n20947 , n14007 , n9779 );
    or g16971 ( n17272 , n4163 , n24973 );
    and g16972 ( n9416 , n3309 , n10536 );
    or g16973 ( n29137 , n28782 , n17030 );
    or g16974 ( n7206 , n8561 , n27865 );
    not g16975 ( n15392 , n17912 );
    or g16976 ( n25085 , n24712 , n27575 );
    not g16977 ( n23868 , n30697 );
    and g16978 ( n9378 , n22134 , n17084 );
    not g16979 ( n12778 , n5679 );
    or g16980 ( n6835 , n5431 , n3857 );
    not g16981 ( n26332 , n30823 );
    not g16982 ( n10835 , n23919 );
    nor g16983 ( n16449 , n6626 , n13425 );
    not g16984 ( n8894 , n9427 );
    not g16985 ( n12128 , n4144 );
    not g16986 ( n13685 , n20955 );
    xnor g16987 ( n1577 , n12880 , n14923 );
    and g16988 ( n9180 , n13071 , n9421 );
    not g16989 ( n24120 , n31287 );
    not g16990 ( n3171 , n13751 );
    and g16991 ( n7977 , n1937 , n10247 );
    not g16992 ( n18619 , n21717 );
    xnor g16993 ( n9517 , n27665 , n17539 );
    and g16994 ( n25594 , n9429 , n25019 );
    and g16995 ( n29098 , n3294 , n19119 );
    xnor g16996 ( n6646 , n2862 , n3432 );
    not g16997 ( n22325 , n28624 );
    xnor g16998 ( n14085 , n13596 , n24008 );
    or g16999 ( n1141 , n2120 , n8164 );
    xnor g17000 ( n23787 , n26613 , n5057 );
    not g17001 ( n24944 , n13196 );
    not g17002 ( n16908 , n13533 );
    xnor g17003 ( n17979 , n25907 , n26262 );
    not g17004 ( n29324 , n25844 );
    not g17005 ( n6436 , n15981 );
    xnor g17006 ( n17945 , n12803 , n3108 );
    not g17007 ( n25872 , n19489 );
    or g17008 ( n18909 , n12427 , n27798 );
    not g17009 ( n30171 , n26713 );
    nor g17010 ( n26383 , n23444 , n2146 );
    xnor g17011 ( n15634 , n25145 , n17342 );
    and g17012 ( n27116 , n19436 , n22899 );
    and g17013 ( n6979 , n7625 , n29938 );
    and g17014 ( n2747 , n1138 , n6675 );
    or g17015 ( n26044 , n15548 , n23178 );
    not g17016 ( n11116 , n27285 );
    xnor g17017 ( n11985 , n13692 , n4562 );
    and g17018 ( n8998 , n8046 , n30365 );
    or g17019 ( n22982 , n22403 , n21573 );
    or g17020 ( n22893 , n16116 , n23691 );
    and g17021 ( n19290 , n9313 , n26249 );
    xnor g17022 ( n5409 , n27908 , n534 );
    and g17023 ( n55 , n1300 , n3669 );
    or g17024 ( n1387 , n24957 , n16742 );
    nor g17025 ( n5367 , n26161 , n29912 );
    xnor g17026 ( n12783 , n6035 , n689 );
    xnor g17027 ( n31165 , n7084 , n17447 );
    nor g17028 ( n15259 , n25040 , n14230 );
    and g17029 ( n16797 , n14528 , n2421 );
    and g17030 ( n30298 , n22955 , n23215 );
    and g17031 ( n29543 , n20806 , n14047 );
    xnor g17032 ( n9857 , n3878 , n17760 );
    not g17033 ( n21757 , n11970 );
    and g17034 ( n22438 , n26282 , n18931 );
    not g17035 ( n3692 , n27885 );
    xnor g17036 ( n7688 , n1177 , n4956 );
    xnor g17037 ( n2185 , n7361 , n19921 );
    not g17038 ( n9478 , n24965 );
    xnor g17039 ( n31350 , n15942 , n26348 );
    or g17040 ( n8047 , n8014 , n13346 );
    xnor g17041 ( n24043 , n31404 , n20553 );
    nor g17042 ( n2037 , n21131 , n3875 );
    or g17043 ( n17045 , n27182 , n29914 );
    or g17044 ( n23575 , n7967 , n17294 );
    and g17045 ( n10660 , n6375 , n10079 );
    not g17046 ( n25869 , n31258 );
    not g17047 ( n16774 , n10635 );
    not g17048 ( n11512 , n18945 );
    or g17049 ( n10182 , n11231 , n29098 );
    and g17050 ( n6898 , n1509 , n18212 );
    xnor g17051 ( n14348 , n17896 , n21386 );
    xnor g17052 ( n23965 , n28877 , n30513 );
    and g17053 ( n5780 , n17140 , n23745 );
    xnor g17054 ( n13003 , n29937 , n9585 );
    or g17055 ( n20745 , n6940 , n18856 );
    and g17056 ( n27875 , n26613 , n23303 );
    or g17057 ( n14275 , n25600 , n26283 );
    and g17058 ( n11277 , n16577 , n19807 );
    not g17059 ( n12401 , n10203 );
    xnor g17060 ( n31258 , n3409 , n23685 );
    xnor g17061 ( n30799 , n27316 , n30808 );
    or g17062 ( n21727 , n29107 , n8322 );
    xnor g17063 ( n8737 , n32022 , n2577 );
    nor g17064 ( n4769 , n20388 , n13554 );
    or g17065 ( n21041 , n6191 , n17835 );
    not g17066 ( n4882 , n24833 );
    nor g17067 ( n17600 , n4821 , n12065 );
    xnor g17068 ( n2987 , n4223 , n11566 );
    xnor g17069 ( n18599 , n24293 , n694 );
    xnor g17070 ( n15890 , n10053 , n13758 );
    xnor g17071 ( n5968 , n6725 , n1366 );
    xnor g17072 ( n17802 , n5506 , n7780 );
    or g17073 ( n25433 , n18730 , n13089 );
    not g17074 ( n22086 , n1934 );
    and g17075 ( n16766 , n1452 , n22705 );
    not g17076 ( n2604 , n25562 );
    not g17077 ( n16261 , n24446 );
    and g17078 ( n28563 , n27931 , n7868 );
    not g17079 ( n1552 , n29390 );
    not g17080 ( n22098 , n4458 );
    not g17081 ( n3013 , n23266 );
    not g17082 ( n29596 , n7943 );
    nor g17083 ( n28391 , n14050 , n5317 );
    and g17084 ( n9660 , n28132 , n31062 );
    xnor g17085 ( n31484 , n6706 , n16124 );
    xnor g17086 ( n3701 , n27007 , n1875 );
    not g17087 ( n29587 , n31711 );
    or g17088 ( n24380 , n24794 , n23173 );
    or g17089 ( n19338 , n6129 , n6182 );
    or g17090 ( n2783 , n25817 , n16857 );
    xnor g17091 ( n32029 , n10020 , n6150 );
    not g17092 ( n30043 , n2834 );
    and g17093 ( n1391 , n14070 , n10955 );
    or g17094 ( n16222 , n10133 , n12724 );
    xnor g17095 ( n18627 , n23004 , n6889 );
    or g17096 ( n2523 , n18082 , n9388 );
    or g17097 ( n31902 , n19419 , n13824 );
    not g17098 ( n10312 , n16139 );
    or g17099 ( n30538 , n18582 , n24905 );
    not g17100 ( n30308 , n3618 );
    not g17101 ( n30948 , n20888 );
    not g17102 ( n16151 , n5531 );
    or g17103 ( n19203 , n28642 , n13155 );
    not g17104 ( n12025 , n21612 );
    xnor g17105 ( n7925 , n26278 , n827 );
    xnor g17106 ( n11613 , n30770 , n18917 );
    xnor g17107 ( n27730 , n16001 , n16321 );
    xnor g17108 ( n6949 , n26640 , n1018 );
    and g17109 ( n26943 , n17011 , n10582 );
    or g17110 ( n27781 , n1499 , n18499 );
    xnor g17111 ( n12223 , n11295 , n29645 );
    xnor g17112 ( n8745 , n12702 , n25936 );
    nor g17113 ( n15185 , n24784 , n18884 );
    xnor g17114 ( n6367 , n30437 , n18209 );
    or g17115 ( n19698 , n3131 , n17641 );
    xnor g17116 ( n5691 , n23029 , n6717 );
    xnor g17117 ( n14638 , n6272 , n21903 );
    xnor g17118 ( n20843 , n1910 , n12018 );
    or g17119 ( n17719 , n13994 , n14733 );
    not g17120 ( n1250 , n6735 );
    xnor g17121 ( n8424 , n18313 , n726 );
    not g17122 ( n3141 , n31023 );
    not g17123 ( n7838 , n11056 );
    or g17124 ( n27604 , n18973 , n31799 );
    xnor g17125 ( n14212 , n23658 , n3831 );
    xnor g17126 ( n5888 , n8429 , n14140 );
    or g17127 ( n24076 , n3599 , n13935 );
    nor g17128 ( n19930 , n17796 , n19534 );
    and g17129 ( n3091 , n25281 , n1004 );
    not g17130 ( n29622 , n158 );
    or g17131 ( n22988 , n3232 , n26076 );
    xnor g17132 ( n31115 , n11607 , n1618 );
    and g17133 ( n1981 , n9248 , n1197 );
    xnor g17134 ( n7687 , n7772 , n11161 );
    not g17135 ( n8586 , n30887 );
    not g17136 ( n17884 , n8232 );
    or g17137 ( n1160 , n3404 , n6824 );
    xnor g17138 ( n17073 , n9335 , n27405 );
    or g17139 ( n29278 , n13711 , n28715 );
    xnor g17140 ( n2074 , n29410 , n24674 );
    not g17141 ( n3968 , n28937 );
    or g17142 ( n24248 , n11957 , n22928 );
    or g17143 ( n16395 , n15270 , n17744 );
    not g17144 ( n17888 , n5800 );
    xnor g17145 ( n27305 , n4369 , n15037 );
    or g17146 ( n18834 , n545 , n17187 );
    or g17147 ( n26543 , n19246 , n10901 );
    or g17148 ( n28073 , n10949 , n9307 );
    xnor g17149 ( n26553 , n30942 , n22224 );
    nor g17150 ( n6732 , n21997 , n18679 );
    not g17151 ( n12692 , n12613 );
    not g17152 ( n18527 , n24490 );
    not g17153 ( n23742 , n879 );
    or g17154 ( n29815 , n18667 , n19632 );
    and g17155 ( n1762 , n28418 , n9196 );
    and g17156 ( n3749 , n20085 , n15754 );
    xnor g17157 ( n30340 , n30645 , n30889 );
    and g17158 ( n19659 , n14621 , n19898 );
    xnor g17159 ( n17138 , n31097 , n22733 );
    not g17160 ( n417 , n11724 );
    or g17161 ( n17659 , n12902 , n10616 );
    not g17162 ( n15176 , n18534 );
    xnor g17163 ( n22936 , n30879 , n19173 );
    xnor g17164 ( n18702 , n21232 , n22149 );
    or g17165 ( n29009 , n12645 , n31865 );
    or g17166 ( n26816 , n21821 , n2827 );
    not g17167 ( n21701 , n23550 );
    or g17168 ( n14294 , n16558 , n2515 );
    or g17169 ( n27468 , n23566 , n7819 );
    not g17170 ( n4383 , n29920 );
    and g17171 ( n18364 , n8587 , n30205 );
    not g17172 ( n30498 , n1002 );
    xnor g17173 ( n1420 , n27093 , n5566 );
    or g17174 ( n30049 , n4795 , n28712 );
    or g17175 ( n14903 , n24209 , n26975 );
    xor g17176 ( n3314 , n9275 , n4418 );
    nor g17177 ( n21462 , n11017 , n8739 );
    or g17178 ( n26426 , n26670 , n19805 );
    or g17179 ( n2307 , n6020 , n968 );
    not g17180 ( n2785 , n12747 );
    not g17181 ( n14787 , n17124 );
    xnor g17182 ( n6709 , n16706 , n31375 );
    and g17183 ( n13872 , n18185 , n28850 );
    not g17184 ( n21165 , n946 );
    and g17185 ( n3947 , n7134 , n27666 );
    or g17186 ( n29127 , n23195 , n9533 );
    not g17187 ( n16736 , n15748 );
    not g17188 ( n16298 , n16706 );
    not g17189 ( n13387 , n9578 );
    not g17190 ( n390 , n31438 );
    and g17191 ( n8038 , n7949 , n26671 );
    or g17192 ( n2249 , n11088 , n8850 );
    or g17193 ( n24052 , n27582 , n21016 );
    xnor g17194 ( n13556 , n15915 , n14977 );
    not g17195 ( n10131 , n27233 );
    or g17196 ( n9440 , n4116 , n28424 );
    xnor g17197 ( n9223 , n6353 , n26483 );
    not g17198 ( n15718 , n27016 );
    not g17199 ( n30967 , n792 );
    xnor g17200 ( n16707 , n8332 , n12500 );
    not g17201 ( n21228 , n8330 );
    not g17202 ( n8155 , n21410 );
    nor g17203 ( n10921 , n13798 , n31583 );
    or g17204 ( n28053 , n1763 , n24417 );
    or g17205 ( n25561 , n4507 , n20819 );
    nor g17206 ( n25659 , n9091 , n31196 );
    not g17207 ( n26924 , n13130 );
    xnor g17208 ( n9173 , n3620 , n11610 );
    not g17209 ( n27578 , n17468 );
    xnor g17210 ( n15183 , n8328 , n16776 );
    nor g17211 ( n2278 , n9239 , n11674 );
    and g17212 ( n31649 , n20587 , n17095 );
    xnor g17213 ( n3008 , n19329 , n14300 );
    xnor g17214 ( n31109 , n29420 , n17334 );
    or g17215 ( n23872 , n26800 , n11042 );
    not g17216 ( n26750 , n8509 );
    not g17217 ( n8514 , n107 );
    not g17218 ( n1639 , n28331 );
    or g17219 ( n17105 , n29100 , n19041 );
    not g17220 ( n16847 , n18002 );
    xnor g17221 ( n31248 , n29342 , n12364 );
    and g17222 ( n30300 , n28114 , n30772 );
    or g17223 ( n9640 , n6340 , n31608 );
    and g17224 ( n20255 , n8829 , n26441 );
    and g17225 ( n8073 , n27324 , n7527 );
    xnor g17226 ( n7094 , n19127 , n981 );
    or g17227 ( n18190 , n13106 , n30888 );
    or g17228 ( n30509 , n7705 , n13454 );
    and g17229 ( n25710 , n26014 , n27044 );
    and g17230 ( n13023 , n11396 , n15680 );
    not g17231 ( n15095 , n31690 );
    not g17232 ( n375 , n142 );
    xnor g17233 ( n4280 , n20920 , n11305 );
    nor g17234 ( n19223 , n22434 , n21316 );
    not g17235 ( n23069 , n26706 );
    xnor g17236 ( n14305 , n22470 , n5113 );
    not g17237 ( n28375 , n25551 );
    or g17238 ( n5460 , n23547 , n31013 );
    not g17239 ( n29746 , n508 );
    not g17240 ( n25064 , n12368 );
    xnor g17241 ( n12317 , n14356 , n2963 );
    and g17242 ( n1763 , n19885 , n12865 );
    and g17243 ( n22056 , n25885 , n30379 );
    not g17244 ( n30131 , n8159 );
    not g17245 ( n14444 , n25999 );
    not g17246 ( n20311 , n12146 );
    not g17247 ( n16972 , n20857 );
    xnor g17248 ( n23925 , n903 , n629 );
    not g17249 ( n886 , n12593 );
    and g17250 ( n13125 , n18631 , n4069 );
    or g17251 ( n9977 , n2982 , n3806 );
    or g17252 ( n11898 , n30669 , n11533 );
    xnor g17253 ( n345 , n22345 , n27805 );
    and g17254 ( n24320 , n14617 , n4275 );
    or g17255 ( n27254 , n4443 , n28182 );
    xnor g17256 ( n21558 , n12823 , n18446 );
    buf g17257 ( n25982 , n11804 );
    and g17258 ( n31213 , n13251 , n1256 );
    or g17259 ( n4558 , n10137 , n8145 );
    and g17260 ( n30654 , n18791 , n3208 );
    xnor g17261 ( n23012 , n19571 , n17863 );
    not g17262 ( n13765 , n26436 );
    xnor g17263 ( n31848 , n29900 , n30320 );
    xnor g17264 ( n8640 , n16969 , n10657 );
    or g17265 ( n6013 , n23133 , n27113 );
    nor g17266 ( n5204 , n561 , n26247 );
    xnor g17267 ( n13950 , n28617 , n7982 );
    not g17268 ( n15356 , n28250 );
    not g17269 ( n9411 , n17969 );
    xnor g17270 ( n3009 , n12319 , n3863 );
    not g17271 ( n23546 , n22665 );
    or g17272 ( n1352 , n17366 , n26074 );
    not g17273 ( n23404 , n805 );
    nor g17274 ( n15950 , n19918 , n24566 );
    not g17275 ( n25092 , n17574 );
    not g17276 ( n22287 , n16586 );
    and g17277 ( n21376 , n3546 , n9793 );
    xnor g17278 ( n23448 , n11498 , n322 );
    not g17279 ( n27366 , n26647 );
    and g17280 ( n25636 , n22420 , n5356 );
    not g17281 ( n9179 , n20236 );
    not g17282 ( n30334 , n3166 );
    not g17283 ( n5411 , n3936 );
    nor g17284 ( n8376 , n19701 , n563 );
    not g17285 ( n15091 , n28872 );
    not g17286 ( n8657 , n25976 );
    xnor g17287 ( n12468 , n17972 , n15858 );
    or g17288 ( n1183 , n27873 , n2282 );
    not g17289 ( n24305 , n11202 );
    or g17290 ( n28838 , n1384 , n6998 );
    xnor g17291 ( n25254 , n14543 , n19274 );
    not g17292 ( n21629 , n1285 );
    xnor g17293 ( n10937 , n28211 , n14489 );
    not g17294 ( n28782 , n18647 );
    or g17295 ( n19151 , n3933 , n6882 );
    and g17296 ( n21987 , n2038 , n31793 );
    not g17297 ( n31926 , n23947 );
    or g17298 ( n1459 , n16441 , n29091 );
    and g17299 ( n22252 , n517 , n3230 );
    xnor g17300 ( n738 , n4739 , n20400 );
    or g17301 ( n7842 , n2187 , n24091 );
    or g17302 ( n3842 , n24158 , n18288 );
    or g17303 ( n10505 , n6429 , n31062 );
    xnor g17304 ( n8222 , n1479 , n3810 );
    not g17305 ( n15687 , n13517 );
    and g17306 ( n13967 , n957 , n19725 );
    buf g17307 ( n20313 , n18995 );
    xnor g17308 ( n8853 , n30917 , n3996 );
    or g17309 ( n1583 , n3444 , n21335 );
    or g17310 ( n13108 , n15402 , n244 );
    and g17311 ( n7750 , n26984 , n5885 );
    and g17312 ( n19749 , n22585 , n8619 );
    nor g17313 ( n31016 , n21264 , n26388 );
    not g17314 ( n1675 , n22429 );
    xnor g17315 ( n23076 , n21910 , n15183 );
    not g17316 ( n13666 , n12187 );
    and g17317 ( n10900 , n29350 , n18571 );
    or g17318 ( n19656 , n10643 , n30426 );
    or g17319 ( n7251 , n7726 , n17097 );
    or g17320 ( n20053 , n11946 , n4858 );
    not g17321 ( n21782 , n5221 );
    nor g17322 ( n28984 , n28417 , n10249 );
    not g17323 ( n30530 , n37 );
    xnor g17324 ( n31348 , n25135 , n22917 );
    xnor g17325 ( n5262 , n28074 , n3976 );
    or g17326 ( n24683 , n13745 , n22220 );
    not g17327 ( n10527 , n21322 );
    not g17328 ( n30013 , n27461 );
    nor g17329 ( n11136 , n9338 , n17739 );
    and g17330 ( n26146 , n23939 , n6668 );
    xnor g17331 ( n25517 , n28517 , n9691 );
    and g17332 ( n28592 , n10652 , n12125 );
    and g17333 ( n29161 , n4938 , n7614 );
    xnor g17334 ( n21467 , n7180 , n21597 );
    not g17335 ( n18450 , n15876 );
    xnor g17336 ( n20071 , n23147 , n14337 );
    not g17337 ( n26856 , n417 );
    nor g17338 ( n18493 , n10490 , n6196 );
    not g17339 ( n25703 , n27267 );
    or g17340 ( n7327 , n18047 , n22993 );
    and g17341 ( n21974 , n23307 , n4971 );
    not g17342 ( n5012 , n13895 );
    or g17343 ( n9384 , n16308 , n22234 );
    not g17344 ( n29298 , n25049 );
    xnor g17345 ( n5220 , n28152 , n23345 );
    not g17346 ( n21443 , n2939 );
    xnor g17347 ( n26224 , n22810 , n22675 );
    and g17348 ( n14692 , n22972 , n7451 );
    and g17349 ( n8885 , n8084 , n14830 );
    and g17350 ( n958 , n20179 , n13584 );
    or g17351 ( n27798 , n5142 , n1429 );
    xnor g17352 ( n28642 , n10135 , n1159 );
    or g17353 ( n19169 , n19211 , n11958 );
    xnor g17354 ( n30119 , n14909 , n4391 );
    or g17355 ( n17050 , n26531 , n17399 );
    nor g17356 ( n8242 , n16746 , n26232 );
    xor g17357 ( n29183 , n13985 , n28397 );
    xnor g17358 ( n12498 , n5453 , n8030 );
    or g17359 ( n3320 , n25455 , n1538 );
    or g17360 ( n1266 , n19142 , n31930 );
    nor g17361 ( n13799 , n17592 , n16142 );
    and g17362 ( n23206 , n30928 , n31169 );
    or g17363 ( n6390 , n24823 , n11563 );
    and g17364 ( n16073 , n2306 , n20948 );
    nor g17365 ( n28479 , n20759 , n28634 );
    xor g17366 ( n10148 , n5526 , n8867 );
    xnor g17367 ( n18401 , n16121 , n10804 );
    not g17368 ( n10786 , n7341 );
    xnor g17369 ( n21429 , n17090 , n31168 );
    xnor g17370 ( n18910 , n30131 , n16516 );
    or g17371 ( n15831 , n15127 , n31702 );
    xnor g17372 ( n14941 , n29035 , n7252 );
    and g17373 ( n30864 , n14075 , n15157 );
    nor g17374 ( n24631 , n9469 , n25291 );
    not g17375 ( n4227 , n28050 );
    or g17376 ( n921 , n17445 , n13516 );
    nor g17377 ( n30341 , n21931 , n14688 );
    xnor g17378 ( n14910 , n9574 , n6422 );
    xnor g17379 ( n13355 , n29079 , n17123 );
    or g17380 ( n20710 , n22095 , n29810 );
    not g17381 ( n31750 , n25414 );
    or g17382 ( n5104 , n15632 , n11545 );
    not g17383 ( n21986 , n14099 );
    not g17384 ( n12147 , n7545 );
    not g17385 ( n19179 , n25577 );
    xnor g17386 ( n23905 , n28006 , n5149 );
    xnor g17387 ( n1353 , n12054 , n1230 );
    not g17388 ( n27972 , n22591 );
    not g17389 ( n4851 , n3964 );
    not g17390 ( n27579 , n13192 );
    or g17391 ( n14644 , n23715 , n5419 );
    not g17392 ( n15130 , n15079 );
    nor g17393 ( n29797 , n5476 , n27466 );
    and g17394 ( n18784 , n14028 , n2611 );
    xor g17395 ( n10555 , n12261 , n14152 );
    xor g17396 ( n170 , n17071 , n7473 );
    or g17397 ( n20984 , n8045 , n6263 );
    xnor g17398 ( n12901 , n14968 , n3548 );
    or g17399 ( n5031 , n7365 , n2182 );
    or g17400 ( n28628 , n29910 , n20508 );
    or g17401 ( n21267 , n9598 , n18426 );
    and g17402 ( n23124 , n21424 , n6295 );
    and g17403 ( n28296 , n27329 , n6268 );
    nor g17404 ( n6301 , n11938 , n11127 );
    xnor g17405 ( n31203 , n22786 , n264 );
    not g17406 ( n29837 , n6223 );
    or g17407 ( n30747 , n10199 , n20302 );
    or g17408 ( n6029 , n12294 , n13076 );
    not g17409 ( n26458 , n22363 );
    xnor g17410 ( n18729 , n5123 , n4052 );
    xnor g17411 ( n13332 , n4269 , n21260 );
    nor g17412 ( n31980 , n8292 , n2690 );
    and g17413 ( n23803 , n12339 , n26426 );
    not g17414 ( n17786 , n22792 );
    not g17415 ( n30944 , n165 );
    and g17416 ( n21823 , n3543 , n28628 );
    or g17417 ( n25041 , n18741 , n13 );
    or g17418 ( n20869 , n30343 , n21266 );
    xnor g17419 ( n3772 , n17203 , n17041 );
    not g17420 ( n26708 , n16997 );
    not g17421 ( n28234 , n19399 );
    xnor g17422 ( n13660 , n6277 , n20645 );
    and g17423 ( n16679 , n23465 , n1885 );
    not g17424 ( n25590 , n10114 );
    or g17425 ( n19589 , n19217 , n9962 );
    xnor g17426 ( n1308 , n20149 , n21749 );
    or g17427 ( n1297 , n18377 , n26509 );
    nor g17428 ( n31086 , n4847 , n9968 );
    and g17429 ( n13066 , n5451 , n30831 );
    not g17430 ( n10351 , n17346 );
    or g17431 ( n23298 , n24733 , n9121 );
    or g17432 ( n27260 , n2744 , n8281 );
    and g17433 ( n19629 , n22330 , n5477 );
    xnor g17434 ( n25551 , n31891 , n12465 );
    not g17435 ( n10655 , n14590 );
    not g17436 ( n8860 , n19220 );
    not g17437 ( n16724 , n27204 );
    or g17438 ( n3712 , n16598 , n28297 );
    not g17439 ( n28942 , n4218 );
    or g17440 ( n19199 , n3688 , n26032 );
    or g17441 ( n22198 , n28142 , n30375 );
    or g17442 ( n1645 , n5488 , n16849 );
    or g17443 ( n16293 , n3070 , n6257 );
    or g17444 ( n12949 , n29934 , n20509 );
    xor g17445 ( n10032 , n13243 , n25926 );
    or g17446 ( n10195 , n16516 , n8159 );
    xnor g17447 ( n23345 , n18119 , n18825 );
    and g17448 ( n17211 , n30407 , n9850 );
    or g17449 ( n30580 , n185 , n8630 );
    xnor g17450 ( n19043 , n30501 , n28300 );
    or g17451 ( n28236 , n16548 , n4083 );
    not g17452 ( n30339 , n21708 );
    or g17453 ( n2897 , n23527 , n14963 );
    xnor g17454 ( n22925 , n2537 , n10939 );
    or g17455 ( n20272 , n7787 , n31708 );
    nor g17456 ( n21004 , n21167 , n10574 );
    not g17457 ( n9263 , n12900 );
    not g17458 ( n7922 , n31755 );
    xnor g17459 ( n1875 , n31571 , n8104 );
    or g17460 ( n23670 , n19400 , n19331 );
    or g17461 ( n3748 , n30067 , n14135 );
    xnor g17462 ( n20042 , n10056 , n28259 );
    and g17463 ( n9419 , n1013 , n6290 );
    xnor g17464 ( n6830 , n6367 , n20556 );
    or g17465 ( n6375 , n26865 , n3941 );
    xnor g17466 ( n11689 , n7210 , n9655 );
    not g17467 ( n7821 , n20485 );
    xnor g17468 ( n26317 , n15193 , n5334 );
    or g17469 ( n15349 , n16815 , n15776 );
    buf g17470 ( n12971 , n14779 );
    not g17471 ( n29841 , n29930 );
    not g17472 ( n19090 , n10125 );
    not g17473 ( n669 , n2570 );
    not g17474 ( n25115 , n3259 );
    not g17475 ( n25766 , n24873 );
    not g17476 ( n7402 , n24649 );
    not g17477 ( n24214 , n3453 );
    not g17478 ( n27267 , n14696 );
    xnor g17479 ( n25367 , n21560 , n27587 );
    and g17480 ( n30721 , n18175 , n801 );
    xnor g17481 ( n19923 , n27306 , n10714 );
    and g17482 ( n26232 , n23569 , n18200 );
    and g17483 ( n19506 , n16138 , n12586 );
    or g17484 ( n4328 , n12694 , n31414 );
    and g17485 ( n13655 , n23146 , n25381 );
    not g17486 ( n21634 , n27964 );
    and g17487 ( n19779 , n11795 , n10320 );
    nor g17488 ( n6176 , n397 , n30486 );
    and g17489 ( n3187 , n3351 , n2471 );
    or g17490 ( n27619 , n11675 , n1612 );
    and g17491 ( n25511 , n5539 , n29025 );
    or g17492 ( n3740 , n29880 , n1949 );
    not g17493 ( n6980 , n19478 );
    or g17494 ( n23451 , n3909 , n31794 );
    xnor g17495 ( n6743 , n7979 , n23994 );
    not g17496 ( n20200 , n31477 );
    not g17497 ( n19100 , n15110 );
    and g17498 ( n9260 , n26107 , n1080 );
    xnor g17499 ( n7031 , n60 , n25299 );
    xnor g17500 ( n29307 , n15054 , n21298 );
    not g17501 ( n9789 , n22836 );
    or g17502 ( n1513 , n13980 , n20714 );
    not g17503 ( n25643 , n22472 );
    xnor g17504 ( n10804 , n3818 , n14206 );
    xnor g17505 ( n27412 , n29584 , n17771 );
    and g17506 ( n2043 , n10428 , n5565 );
    not g17507 ( n19581 , n7151 );
    xor g17508 ( n15222 , n29903 , n16310 );
    and g17509 ( n10756 , n31598 , n29256 );
    nor g17510 ( n12567 , n21953 , n22372 );
    not g17511 ( n12813 , n5560 );
    not g17512 ( n5610 , n20253 );
    xnor g17513 ( n20205 , n22332 , n23335 );
    xnor g17514 ( n26461 , n24116 , n8104 );
    and g17515 ( n28425 , n18549 , n3345 );
    xor g17516 ( n27196 , n15230 , n5783 );
    or g17517 ( n2619 , n14751 , n28629 );
    not g17518 ( n22145 , n3173 );
    xnor g17519 ( n1021 , n28433 , n14035 );
    and g17520 ( n4486 , n15773 , n15503 );
    or g17521 ( n6887 , n27039 , n746 );
    and g17522 ( n3200 , n29748 , n2427 );
    not g17523 ( n30088 , n16609 );
    or g17524 ( n16748 , n29249 , n3588 );
    xnor g17525 ( n23824 , n16828 , n20180 );
    or g17526 ( n12249 , n19464 , n2799 );
    nor g17527 ( n16015 , n20789 , n5221 );
    not g17528 ( n14995 , n24463 );
    not g17529 ( n13771 , n19710 );
    and g17530 ( n10240 , n8484 , n3312 );
    not g17531 ( n9976 , n4711 );
    and g17532 ( n2932 , n23816 , n18129 );
    nor g17533 ( n280 , n20269 , n21229 );
    xnor g17534 ( n4606 , n26936 , n30285 );
    or g17535 ( n21630 , n29912 , n8510 );
    xnor g17536 ( n16911 , n4117 , n20967 );
    or g17537 ( n234 , n11984 , n4425 );
    xnor g17538 ( n20446 , n6415 , n3106 );
    xnor g17539 ( n11947 , n15685 , n12497 );
    nor g17540 ( n26043 , n27602 , n23828 );
    and g17541 ( n29419 , n17874 , n25769 );
    nor g17542 ( n23791 , n29391 , n12418 );
    not g17543 ( n4883 , n21940 );
    not g17544 ( n31951 , n5273 );
    xnor g17545 ( n16170 , n17486 , n6880 );
    xnor g17546 ( n22695 , n23205 , n20357 );
    xor g17547 ( n30697 , n15160 , n11994 );
    not g17548 ( n19897 , n26545 );
    and g17549 ( n28235 , n10821 , n12761 );
    xnor g17550 ( n25173 , n1924 , n31298 );
    not g17551 ( n12427 , n13897 );
    or g17552 ( n31658 , n30831 , n28770 );
    xnor g17553 ( n23388 , n25621 , n11850 );
    xnor g17554 ( n30962 , n9310 , n10737 );
    xnor g17555 ( n8314 , n22109 , n23032 );
    not g17556 ( n26705 , n27534 );
    and g17557 ( n28055 , n5526 , n8867 );
    or g17558 ( n14476 , n3189 , n19315 );
    not g17559 ( n20572 , n29918 );
    xnor g17560 ( n6680 , n27831 , n7412 );
    not g17561 ( n18339 , n22645 );
    or g17562 ( n19052 , n18376 , n18194 );
    and g17563 ( n16827 , n4965 , n31925 );
    xnor g17564 ( n14817 , n49 , n20866 );
    xnor g17565 ( n21377 , n10392 , n7037 );
    nor g17566 ( n11124 , n26403 , n14238 );
    not g17567 ( n14537 , n27805 );
    and g17568 ( n7917 , n17581 , n79 );
    or g17569 ( n15615 , n19740 , n2239 );
    xnor g17570 ( n8379 , n15752 , n4993 );
    not g17571 ( n11781 , n21131 );
    xnor g17572 ( n2548 , n9262 , n9818 );
    and g17573 ( n20646 , n27001 , n8575 );
    or g17574 ( n6022 , n17157 , n19552 );
    not g17575 ( n18096 , n13924 );
    xnor g17576 ( n14930 , n21774 , n17416 );
    and g17577 ( n4860 , n30190 , n3318 );
    xnor g17578 ( n30892 , n9631 , n20937 );
    not g17579 ( n25452 , n16815 );
    xnor g17580 ( n13308 , n29161 , n22342 );
    nor g17581 ( n23078 , n3442 , n15888 );
    not g17582 ( n23178 , n2772 );
    or g17583 ( n14419 , n11051 , n383 );
    or g17584 ( n27051 , n16933 , n10861 );
    not g17585 ( n29770 , n16862 );
    not g17586 ( n8029 , n4554 );
    or g17587 ( n15725 , n9889 , n22924 );
    xnor g17588 ( n22123 , n9272 , n17250 );
    xnor g17589 ( n26891 , n9611 , n27546 );
    not g17590 ( n1440 , n12926 );
    or g17591 ( n23147 , n30883 , n13848 );
    nor g17592 ( n28981 , n29569 , n2660 );
    not g17593 ( n31708 , n9145 );
    or g17594 ( n10579 , n8104 , n5986 );
    not g17595 ( n5827 , n23926 );
    xnor g17596 ( n2995 , n15276 , n21405 );
    xnor g17597 ( n1120 , n22488 , n8811 );
    and g17598 ( n7704 , n27042 , n10326 );
    nor g17599 ( n4116 , n26536 , n19593 );
    and g17600 ( n22409 , n10167 , n25184 );
    not g17601 ( n15108 , n28433 );
    xnor g17602 ( n5817 , n10405 , n5273 );
    xnor g17603 ( n1524 , n23222 , n28625 );
    or g17604 ( n19906 , n14859 , n22780 );
    not g17605 ( n9325 , n22295 );
    not g17606 ( n10492 , n4397 );
    and g17607 ( n9546 , n27603 , n5624 );
    and g17608 ( n837 , n25887 , n4424 );
    or g17609 ( n22651 , n22632 , n6358 );
    xnor g17610 ( n13325 , n4603 , n13925 );
    xnor g17611 ( n10485 , n31075 , n28178 );
    xnor g17612 ( n16091 , n4948 , n17489 );
    xnor g17613 ( n25164 , n5803 , n6838 );
    nor g17614 ( n26205 , n24910 , n10812 );
    not g17615 ( n3933 , n16075 );
    not g17616 ( n2212 , n25189 );
    not g17617 ( n17748 , n17601 );
    and g17618 ( n16017 , n18711 , n17624 );
    xnor g17619 ( n11931 , n2379 , n4590 );
    not g17620 ( n13532 , n16615 );
    xnor g17621 ( n20556 , n14429 , n25419 );
    not g17622 ( n17407 , n10411 );
    not g17623 ( n4583 , n4213 );
    or g17624 ( n15978 , n28169 , n17426 );
    or g17625 ( n1224 , n936 , n653 );
    and g17626 ( n6164 , n19403 , n31052 );
    nor g17627 ( n20368 , n31957 , n3727 );
    not g17628 ( n21321 , n9279 );
    xnor g17629 ( n16579 , n13454 , n8014 );
    nor g17630 ( n19439 , n18764 , n30866 );
    xnor g17631 ( n10358 , n22565 , n29448 );
    or g17632 ( n29657 , n17617 , n7542 );
    not g17633 ( n23474 , n8918 );
    not g17634 ( n935 , n16523 );
    or g17635 ( n18931 , n21316 , n24255 );
    xnor g17636 ( n17640 , n15194 , n25123 );
    or g17637 ( n26679 , n5988 , n25588 );
    xnor g17638 ( n16703 , n22313 , n28024 );
    buf g17639 ( n8133 , n28827 );
    xnor g17640 ( n21007 , n2900 , n19621 );
    not g17641 ( n21379 , n26312 );
    not g17642 ( n2183 , n29441 );
    xnor g17643 ( n27315 , n5398 , n15890 );
    not g17644 ( n25587 , n10490 );
    xnor g17645 ( n13612 , n14447 , n29867 );
    and g17646 ( n7818 , n18009 , n14639 );
    or g17647 ( n15765 , n14352 , n30027 );
    not g17648 ( n28532 , n25493 );
    xnor g17649 ( n24689 , n21439 , n20011 );
    and g17650 ( n27311 , n28987 , n5131 );
    xnor g17651 ( n20199 , n12710 , n7459 );
    not g17652 ( n451 , n5948 );
    or g17653 ( n11357 , n28420 , n30767 );
    xnor g17654 ( n31199 , n519 , n16131 );
    not g17655 ( n24961 , n5086 );
    xnor g17656 ( n12260 , n18193 , n11979 );
    and g17657 ( n3060 , n12875 , n7372 );
    xnor g17658 ( n9723 , n832 , n15785 );
    or g17659 ( n28747 , n218 , n31887 );
    nor g17660 ( n28328 , n9892 , n18286 );
    nor g17661 ( n5331 , n20815 , n13643 );
    not g17662 ( n25488 , n22598 );
    and g17663 ( n22933 , n32008 , n14663 );
    xnor g17664 ( n803 , n715 , n13906 );
    or g17665 ( n9779 , n20043 , n31205 );
    not g17666 ( n368 , n1707 );
    not g17667 ( n17930 , n3854 );
    nor g17668 ( n8313 , n26256 , n3283 );
    not g17669 ( n26409 , n1497 );
    or g17670 ( n23881 , n23581 , n14462 );
    and g17671 ( n6583 , n5284 , n2547 );
    or g17672 ( n9815 , n16475 , n17344 );
    nor g17673 ( n1608 , n28486 , n6097 );
    not g17674 ( n11064 , n23024 );
    and g17675 ( n10207 , n29321 , n5752 );
    and g17676 ( n16605 , n14736 , n26519 );
    not g17677 ( n19228 , n29761 );
    or g17678 ( n2012 , n14579 , n4714 );
    not g17679 ( n21647 , n1109 );
    and g17680 ( n23993 , n4867 , n3493 );
    or g17681 ( n11699 , n9224 , n12470 );
    not g17682 ( n8265 , n11619 );
    xnor g17683 ( n17853 , n21934 , n10327 );
    not g17684 ( n5293 , n10647 );
    or g17685 ( n3414 , n24435 , n16465 );
    xnor g17686 ( n29522 , n8597 , n13352 );
    or g17687 ( n14043 , n12189 , n2154 );
    not g17688 ( n31739 , n18227 );
    and g17689 ( n28324 , n29844 , n17757 );
    or g17690 ( n17673 , n11505 , n5608 );
    not g17691 ( n22049 , n15458 );
    xnor g17692 ( n28847 , n6306 , n10477 );
    not g17693 ( n10102 , n24970 );
    xnor g17694 ( n1791 , n6331 , n8321 );
    nor g17695 ( n28511 , n11745 , n29061 );
    and g17696 ( n20425 , n1627 , n19122 );
    not g17697 ( n4446 , n15433 );
    or g17698 ( n29227 , n29164 , n25349 );
    and g17699 ( n6999 , n1853 , n10949 );
    and g17700 ( n7595 , n25754 , n19868 );
    and g17701 ( n15752 , n22117 , n633 );
    not g17702 ( n3471 , n15710 );
    not g17703 ( n622 , n26444 );
    nor g17704 ( n23157 , n19125 , n20156 );
    xnor g17705 ( n14065 , n16080 , n11771 );
    not g17706 ( n30921 , n29462 );
    not g17707 ( n14931 , n1856 );
    or g17708 ( n16473 , n2713 , n715 );
    not g17709 ( n14266 , n19516 );
    xnor g17710 ( n7104 , n11819 , n4659 );
    not g17711 ( n25562 , n28066 );
    not g17712 ( n9021 , n13980 );
    nor g17713 ( n6378 , n28828 , n31070 );
    or g17714 ( n1221 , n3036 , n13017 );
    not g17715 ( n16386 , n27569 );
    xnor g17716 ( n3419 , n5479 , n27761 );
    not g17717 ( n5699 , n2048 );
    and g17718 ( n20586 , n26010 , n5423 );
    buf g17719 ( n11584 , n28531 );
    not g17720 ( n9508 , n22369 );
    and g17721 ( n23279 , n11188 , n4183 );
    not g17722 ( n27554 , n2968 );
    or g17723 ( n4962 , n10139 , n25760 );
    xnor g17724 ( n5135 , n886 , n10356 );
    and g17725 ( n1383 , n31132 , n8560 );
    and g17726 ( n27146 , n21802 , n25830 );
    or g17727 ( n11941 , n7333 , n29835 );
    xnor g17728 ( n24019 , n1020 , n12210 );
    xor g17729 ( n21728 , n1327 , n12998 );
    or g17730 ( n8435 , n26786 , n17970 );
    and g17731 ( n11216 , n29334 , n14921 );
    or g17732 ( n30205 , n2683 , n17506 );
    not g17733 ( n23103 , n11767 );
    and g17734 ( n4535 , n27891 , n25981 );
    not g17735 ( n24435 , n23886 );
    or g17736 ( n21366 , n11921 , n7026 );
    not g17737 ( n22606 , n8354 );
    and g17738 ( n11487 , n25835 , n8993 );
    and g17739 ( n10399 , n1586 , n13392 );
    or g17740 ( n3198 , n19035 , n31734 );
    not g17741 ( n16041 , n11121 );
    xnor g17742 ( n28978 , n28285 , n7188 );
    not g17743 ( n19093 , n30785 );
    and g17744 ( n17447 , n26384 , n15697 );
    xnor g17745 ( n3265 , n5483 , n763 );
    not g17746 ( n23274 , n24243 );
    not g17747 ( n4249 , n18920 );
    or g17748 ( n18607 , n15146 , n31947 );
    not g17749 ( n26481 , n5275 );
    xnor g17750 ( n23326 , n12387 , n1921 );
    nor g17751 ( n31046 , n25288 , n17965 );
    or g17752 ( n31795 , n31509 , n22024 );
    not g17753 ( n11572 , n22021 );
    or g17754 ( n23242 , n27655 , n21878 );
    not g17755 ( n11943 , n29330 );
    and g17756 ( n4699 , n31480 , n21366 );
    xnor g17757 ( n26012 , n2717 , n12712 );
    nor g17758 ( n3302 , n21228 , n30629 );
    or g17759 ( n23933 , n24331 , n2251 );
    or g17760 ( n19636 , n5281 , n10734 );
    xnor g17761 ( n10377 , n18361 , n3080 );
    and g17762 ( n3662 , n23682 , n12589 );
    xnor g17763 ( n21014 , n29336 , n5113 );
    not g17764 ( n20177 , n13640 );
    or g17765 ( n15918 , n6250 , n646 );
    not g17766 ( n2076 , n18633 );
    not g17767 ( n22079 , n31787 );
    and g17768 ( n14752 , n15834 , n1225 );
    xnor g17769 ( n6106 , n28009 , n21594 );
    or g17770 ( n20037 , n11034 , n13474 );
    xnor g17771 ( n29184 , n9143 , n17224 );
    not g17772 ( n18117 , n4650 );
    and g17773 ( n31471 , n17104 , n4274 );
    xnor g17774 ( n27193 , n23040 , n2939 );
    xnor g17775 ( n29322 , n19044 , n28894 );
    xnor g17776 ( n6705 , n27152 , n26343 );
    not g17777 ( n9482 , n8252 );
    or g17778 ( n29250 , n10981 , n6551 );
    not g17779 ( n21482 , n27002 );
    or g17780 ( n22613 , n17291 , n14195 );
    and g17781 ( n16268 , n20990 , n30429 );
    xnor g17782 ( n9563 , n5000 , n16043 );
    nor g17783 ( n24661 , n15204 , n29596 );
    or g17784 ( n8551 , n4098 , n27340 );
    and g17785 ( n27060 , n27332 , n14846 );
    or g17786 ( n16762 , n11124 , n11371 );
    or g17787 ( n15423 , n9846 , n21740 );
    nor g17788 ( n973 , n24486 , n25289 );
    nor g17789 ( n7607 , n25246 , n22861 );
    nor g17790 ( n19957 , n3563 , n5866 );
    or g17791 ( n7393 , n24196 , n12969 );
    xnor g17792 ( n20954 , n20179 , n20237 );
    or g17793 ( n11731 , n10981 , n3854 );
    not g17794 ( n18919 , n28756 );
    or g17795 ( n31364 , n30204 , n26305 );
    xnor g17796 ( n17285 , n5946 , n26602 );
    and g17797 ( n696 , n26681 , n26907 );
    or g17798 ( n30993 , n7382 , n13178 );
    xnor g17799 ( n30026 , n7619 , n12625 );
    buf g17800 ( n13318 , n29073 );
    not g17801 ( n30409 , n21911 );
    and g17802 ( n27303 , n4618 , n9509 );
    or g17803 ( n26520 , n10554 , n13757 );
    and g17804 ( n17662 , n22263 , n23711 );
    not g17805 ( n28117 , n11303 );
    nor g17806 ( n5134 , n31940 , n22792 );
    xnor g17807 ( n13184 , n1013 , n26678 );
    or g17808 ( n19320 , n11264 , n9782 );
    or g17809 ( n22162 , n29460 , n26016 );
    and g17810 ( n11864 , n27394 , n4688 );
    not g17811 ( n12118 , n17651 );
    or g17812 ( n24511 , n29307 , n4503 );
    xnor g17813 ( n26268 , n17228 , n4127 );
    or g17814 ( n14459 , n7586 , n30508 );
    xnor g17815 ( n6809 , n16989 , n15574 );
    xnor g17816 ( n13164 , n29596 , n7184 );
    not g17817 ( n25747 , n29830 );
    not g17818 ( n22774 , n5951 );
    and g17819 ( n22685 , n5220 , n10474 );
    nor g17820 ( n26019 , n22806 , n4240 );
    xnor g17821 ( n30320 , n6872 , n3267 );
    or g17822 ( n9337 , n18730 , n1864 );
    and g17823 ( n11607 , n17792 , n19993 );
    nor g17824 ( n16197 , n18955 , n4498 );
    and g17825 ( n9438 , n7633 , n9459 );
    or g17826 ( n24878 , n13941 , n20369 );
    xnor g17827 ( n814 , n13258 , n15774 );
    xnor g17828 ( n26130 , n20628 , n22346 );
    nor g17829 ( n8177 , n23289 , n9035 );
    not g17830 ( n12775 , n1154 );
    not g17831 ( n23893 , n3312 );
    or g17832 ( n15696 , n14526 , n8984 );
    xnor g17833 ( n30469 , n97 , n2150 );
    nor g17834 ( n5292 , n21404 , n4464 );
    or g17835 ( n25969 , n28408 , n29171 );
    and g17836 ( n20229 , n1955 , n12179 );
    xnor g17837 ( n22346 , n11462 , n2862 );
    xnor g17838 ( n27152 , n22872 , n30506 );
    not g17839 ( n13724 , n25760 );
    xnor g17840 ( n30010 , n31446 , n19538 );
    not g17841 ( n1853 , n13833 );
    and g17842 ( n3279 , n5522 , n8982 );
    or g17843 ( n29492 , n28950 , n16833 );
    xnor g17844 ( n22256 , n27479 , n9481 );
    xnor g17845 ( n8617 , n1518 , n10676 );
    xnor g17846 ( n10544 , n6108 , n11512 );
    not g17847 ( n6437 , n553 );
    and g17848 ( n16955 , n25922 , n20979 );
    xnor g17849 ( n14666 , n20488 , n23941 );
    or g17850 ( n5740 , n21329 , n16179 );
    xnor g17851 ( n31579 , n30560 , n6097 );
    not g17852 ( n657 , n1856 );
    or g17853 ( n25009 , n14287 , n13560 );
    or g17854 ( n16217 , n15436 , n29218 );
    and g17855 ( n7537 , n3236 , n7486 );
    not g17856 ( n11869 , n21132 );
    xnor g17857 ( n19882 , n14128 , n25809 );
    or g17858 ( n3358 , n657 , n12489 );
    and g17859 ( n24157 , n24399 , n14644 );
    xnor g17860 ( n20384 , n5312 , n9482 );
    not g17861 ( n2438 , n14841 );
    nor g17862 ( n15312 , n19839 , n29812 );
    and g17863 ( n22458 , n4885 , n11330 );
    not g17864 ( n16122 , n12849 );
    and g17865 ( n10855 , n12829 , n2701 );
    xnor g17866 ( n1132 , n18935 , n19858 );
    not g17867 ( n24276 , n2010 );
    or g17868 ( n26928 , n1337 , n8609 );
    and g17869 ( n27649 , n31425 , n12871 );
    and g17870 ( n4969 , n26141 , n9833 );
    not g17871 ( n9635 , n12856 );
    or g17872 ( n7685 , n24298 , n20439 );
    not g17873 ( n31966 , n13735 );
    xnor g17874 ( n17916 , n28740 , n15372 );
    and g17875 ( n3537 , n19640 , n8395 );
    or g17876 ( n26133 , n28022 , n10890 );
    not g17877 ( n1439 , n20069 );
    or g17878 ( n29077 , n14011 , n2871 );
    not g17879 ( n5028 , n5652 );
    and g17880 ( n4121 , n2391 , n2637 );
    xnor g17881 ( n17894 , n27218 , n18760 );
    and g17882 ( n5172 , n4999 , n10504 );
    or g17883 ( n26058 , n25485 , n15168 );
    nor g17884 ( n4224 , n899 , n8491 );
    and g17885 ( n20223 , n3699 , n29769 );
    or g17886 ( n23583 , n22750 , n26949 );
    or g17887 ( n3513 , n11793 , n31621 );
    not g17888 ( n17950 , n8200 );
    nor g17889 ( n7081 , n10949 , n3501 );
    or g17890 ( n343 , n26019 , n1780 );
    xnor g17891 ( n25691 , n16181 , n19228 );
    not g17892 ( n17684 , n5007 );
    xnor g17893 ( n13399 , n9194 , n28640 );
    not g17894 ( n20575 , n13492 );
    or g17895 ( n13874 , n10216 , n22387 );
    not g17896 ( n19905 , n19200 );
    and g17897 ( n23467 , n8527 , n6747 );
    xnor g17898 ( n5742 , n13879 , n15586 );
    or g17899 ( n9082 , n31369 , n25857 );
    nor g17900 ( n9702 , n20854 , n9345 );
    xnor g17901 ( n9555 , n21261 , n21963 );
    nor g17902 ( n14284 , n30972 , n1266 );
    not g17903 ( n27309 , n299 );
    and g17904 ( n16996 , n12984 , n30110 );
    not g17905 ( n18398 , n3280 );
    xnor g17906 ( n24621 , n24046 , n7701 );
    not g17907 ( n31875 , n27818 );
    nor g17908 ( n2498 , n3810 , n4847 );
    and g17909 ( n19305 , n25317 , n2493 );
    xnor g17910 ( n9864 , n29715 , n12320 );
    xnor g17911 ( n23775 , n25717 , n27694 );
    not g17912 ( n25974 , n10357 );
    and g17913 ( n19599 , n18074 , n23984 );
    or g17914 ( n14608 , n18498 , n8354 );
    and g17915 ( n7240 , n10564 , n2869 );
    or g17916 ( n4186 , n25590 , n20955 );
    or g17917 ( n28206 , n10546 , n4809 );
    not g17918 ( n4220 , n20764 );
    or g17919 ( n25875 , n27266 , n222 );
    nor g17920 ( n8293 , n12025 , n2386 );
    nor g17921 ( n26734 , n5018 , n29157 );
    xnor g17922 ( n20613 , n13315 , n24784 );
    or g17923 ( n17922 , n18008 , n6333 );
    and g17924 ( n28033 , n30091 , n9081 );
    not g17925 ( n30994 , n27381 );
    not g17926 ( n736 , n2920 );
    buf g17927 ( n14373 , n18623 );
    not g17928 ( n16045 , n15125 );
    or g17929 ( n20298 , n28915 , n18694 );
    or g17930 ( n27864 , n18714 , n1087 );
    xnor g17931 ( n29981 , n16624 , n30772 );
    not g17932 ( n23914 , n25721 );
    nor g17933 ( n29133 , n24132 , n21044 );
    xnor g17934 ( n26329 , n12668 , n26894 );
    not g17935 ( n18557 , n22970 );
    and g17936 ( n25948 , n21814 , n30936 );
    xnor g17937 ( n3393 , n2740 , n30541 );
    or g17938 ( n17092 , n28653 , n12884 );
    and g17939 ( n31485 , n22964 , n9539 );
    and g17940 ( n21884 , n10874 , n10314 );
    xnor g17941 ( n18644 , n5392 , n5020 );
    xnor g17942 ( n18662 , n16797 , n4652 );
    or g17943 ( n5829 , n25940 , n11902 );
    xnor g17944 ( n15839 , n2939 , n27534 );
    or g17945 ( n1402 , n18771 , n18767 );
    not g17946 ( n21386 , n12122 );
    and g17947 ( n13218 , n16561 , n2135 );
    xnor g17948 ( n15105 , n26601 , n23046 );
    or g17949 ( n28263 , n2925 , n23659 );
    or g17950 ( n11447 , n18396 , n14730 );
    xnor g17951 ( n21889 , n28121 , n29764 );
    xnor g17952 ( n13075 , n5835 , n8900 );
    xnor g17953 ( n10353 , n11748 , n29494 );
    and g17954 ( n10018 , n6364 , n1639 );
    or g17955 ( n27600 , n30956 , n22971 );
    xor g17956 ( n587 , n8471 , n24006 );
    xnor g17957 ( n6939 , n10946 , n29615 );
    not g17958 ( n10013 , n30794 );
    or g17959 ( n20423 , n27279 , n27137 );
    xnor g17960 ( n12385 , n8034 , n23741 );
    and g17961 ( n6077 , n10401 , n11536 );
    not g17962 ( n23001 , n24336 );
    or g17963 ( n13208 , n31919 , n12945 );
    not g17964 ( n23276 , n13729 );
    xnor g17965 ( n28432 , n28787 , n17468 );
    not g17966 ( n26745 , n138 );
    not g17967 ( n19262 , n6056 );
    not g17968 ( n29440 , n25548 );
    xnor g17969 ( n30279 , n25935 , n3570 );
    xnor g17970 ( n23164 , n19954 , n20900 );
    xor g17971 ( n15521 , n27005 , n20459 );
    or g17972 ( n24215 , n19490 , n25120 );
    not g17973 ( n14720 , n11327 );
    not g17974 ( n21350 , n28431 );
    nor g17975 ( n12172 , n10363 , n4525 );
    or g17976 ( n31282 , n12328 , n29110 );
    or g17977 ( n23994 , n14183 , n19488 );
    not g17978 ( n2176 , n5149 );
    nor g17979 ( n4873 , n11153 , n24585 );
    and g17980 ( n14452 , n12221 , n30275 );
    and g17981 ( n24973 , n783 , n13593 );
    and g17982 ( n11620 , n21405 , n31131 );
    xnor g17983 ( n2703 , n9226 , n31057 );
    not g17984 ( n4582 , n9948 );
    or g17985 ( n8498 , n3691 , n14475 );
    xnor g17986 ( n1429 , n16397 , n6797 );
    not g17987 ( n20113 , n19183 );
    nor g17988 ( n13538 , n28644 , n6109 );
    and g17989 ( n16533 , n14567 , n19279 );
    not g17990 ( n4821 , n24415 );
    not g17991 ( n5773 , n25828 );
    or g17992 ( n15403 , n21583 , n2786 );
    nor g17993 ( n1403 , n27737 , n23649 );
    or g17994 ( n17535 , n11925 , n5615 );
    xnor g17995 ( n11592 , n21661 , n24289 );
    or g17996 ( n5557 , n24788 , n29008 );
    nor g17997 ( n682 , n22809 , n28729 );
    xnor g17998 ( n6574 , n23862 , n8278 );
    not g17999 ( n19655 , n4779 );
    or g18000 ( n31564 , n16034 , n31680 );
    or g18001 ( n16614 , n21999 , n13913 );
    not g18002 ( n3119 , n10229 );
    and g18003 ( n4785 , n4094 , n13965 );
    or g18004 ( n28980 , n19355 , n11312 );
    xnor g18005 ( n14821 , n8730 , n11565 );
    not g18006 ( n15813 , n24363 );
    not g18007 ( n8341 , n11149 );
    xnor g18008 ( n4349 , n17183 , n12364 );
    not g18009 ( n16910 , n23539 );
    nor g18010 ( n18011 , n8686 , n9396 );
    and g18011 ( n28323 , n14755 , n14030 );
    and g18012 ( n16812 , n26563 , n17645 );
    nor g18013 ( n5614 , n7314 , n28264 );
    xnor g18014 ( n21684 , n9823 , n22940 );
    and g18015 ( n18309 , n9614 , n13445 );
    or g18016 ( n5863 , n18957 , n12521 );
    xnor g18017 ( n23441 , n5827 , n29145 );
    or g18018 ( n15702 , n29119 , n5194 );
    not g18019 ( n13510 , n18391 );
    xor g18020 ( n28988 , n18752 , n8733 );
    nor g18021 ( n428 , n8479 , n10682 );
    nor g18022 ( n17543 , n6306 , n11375 );
    xnor g18023 ( n31447 , n16913 , n21320 );
    and g18024 ( n23525 , n18066 , n13691 );
    nor g18025 ( n13860 , n31462 , n5715 );
    or g18026 ( n1245 , n9069 , n21079 );
    xnor g18027 ( n6236 , n7919 , n20969 );
    or g18028 ( n2504 , n18076 , n13605 );
    not g18029 ( n13563 , n10943 );
    not g18030 ( n29827 , n16763 );
    or g18031 ( n15313 , n27221 , n8479 );
    or g18032 ( n29167 , n24130 , n6924 );
    xnor g18033 ( n15274 , n10136 , n17832 );
    and g18034 ( n24933 , n25270 , n24847 );
    xnor g18035 ( n21862 , n29183 , n5801 );
    or g18036 ( n8417 , n30595 , n11198 );
    not g18037 ( n25970 , n7799 );
    not g18038 ( n1307 , n3046 );
    nor g18039 ( n15700 , n10521 , n25089 );
    buf g18040 ( n5895 , n16288 );
    not g18041 ( n27440 , n31881 );
    not g18042 ( n14523 , n18389 );
    or g18043 ( n7994 , n2356 , n26767 );
    xnor g18044 ( n13546 , n7083 , n16200 );
    and g18045 ( n30082 , n19713 , n11013 );
    not g18046 ( n14577 , n15396 );
    or g18047 ( n8280 , n22177 , n3050 );
    not g18048 ( n20692 , n3047 );
    or g18049 ( n6728 , n14992 , n14648 );
    and g18050 ( n26451 , n11106 , n20528 );
    and g18051 ( n7156 , n22721 , n2876 );
    or g18052 ( n564 , n11574 , n1524 );
    not g18053 ( n28088 , n9183 );
    and g18054 ( n29962 , n30671 , n10744 );
    or g18055 ( n19014 , n10268 , n14731 );
    not g18056 ( n31140 , n7968 );
    or g18057 ( n1925 , n5281 , n24003 );
    xnor g18058 ( n22856 , n29789 , n19797 );
    not g18059 ( n3563 , n4187 );
    not g18060 ( n4658 , n16308 );
    nor g18061 ( n12050 , n20452 , n12717 );
    xnor g18062 ( n5071 , n2566 , n11262 );
    xnor g18063 ( n548 , n12998 , n7473 );
    or g18064 ( n6382 , n31782 , n17842 );
    xnor g18065 ( n1587 , n27256 , n30231 );
    xnor g18066 ( n14906 , n1845 , n9311 );
    or g18067 ( n1357 , n23744 , n9328 );
    not g18068 ( n14634 , n15298 );
    not g18069 ( n5953 , n22529 );
    not g18070 ( n13388 , n6165 );
    or g18071 ( n18215 , n31559 , n11569 );
    xnor g18072 ( n3023 , n30045 , n6422 );
    nor g18073 ( n26564 , n23964 , n27946 );
    or g18074 ( n6606 , n29293 , n25720 );
    nor g18075 ( n5039 , n14014 , n6952 );
    or g18076 ( n14626 , n5811 , n10240 );
    xnor g18077 ( n31741 , n17721 , n28272 );
    or g18078 ( n11431 , n16231 , n19613 );
    xor g18079 ( n1507 , n30912 , n23299 );
    and g18080 ( n5389 , n19568 , n16896 );
    or g18081 ( n27507 , n16856 , n154 );
    xnor g18082 ( n2809 , n9429 , n20196 );
    or g18083 ( n31738 , n5917 , n6087 );
    not g18084 ( n20225 , n7444 );
    xnor g18085 ( n4238 , n28317 , n26819 );
    not g18086 ( n3175 , n18027 );
    xor g18087 ( n24703 , n16814 , n10320 );
    or g18088 ( n19715 , n575 , n29794 );
    or g18089 ( n15208 , n27322 , n4082 );
    or g18090 ( n10174 , n21317 , n10662 );
    not g18091 ( n31728 , n15460 );
    nor g18092 ( n12166 , n1206 , n20830 );
    xnor g18093 ( n9975 , n17217 , n24018 );
    not g18094 ( n528 , n26433 );
    xnor g18095 ( n4579 , n21886 , n19352 );
    not g18096 ( n28230 , n31460 );
    not g18097 ( n12935 , n7539 );
    xor g18098 ( n15863 , n11032 , n27409 );
    xnor g18099 ( n28367 , n1125 , n7637 );
    nor g18100 ( n3771 , n29764 , n10243 );
    and g18101 ( n19097 , n24143 , n10454 );
    or g18102 ( n4734 , n5320 , n24261 );
    and g18103 ( n28427 , n28919 , n19102 );
    xnor g18104 ( n189 , n30597 , n26670 );
    xnor g18105 ( n23435 , n21116 , n19701 );
    and g18106 ( n24007 , n29704 , n5214 );
    not g18107 ( n3603 , n16910 );
    or g18108 ( n14891 , n23681 , n23456 );
    xnor g18109 ( n21282 , n27692 , n11252 );
    xnor g18110 ( n16338 , n1872 , n8126 );
    xnor g18111 ( n15369 , n26131 , n31095 );
    nor g18112 ( n23955 , n18058 , n16280 );
    and g18113 ( n23222 , n24123 , n23746 );
    and g18114 ( n14412 , n7556 , n628 );
    and g18115 ( n8729 , n20423 , n23105 );
    xnor g18116 ( n23540 , n6644 , n8627 );
    xnor g18117 ( n13360 , n11652 , n31831 );
    nor g18118 ( n2093 , n14872 , n6123 );
    not g18119 ( n13802 , n15738 );
    xnor g18120 ( n18810 , n19204 , n15421 );
    or g18121 ( n28377 , n24523 , n3458 );
    xnor g18122 ( n23978 , n23333 , n2663 );
    not g18123 ( n1350 , n4579 );
    not g18124 ( n12202 , n23633 );
    not g18125 ( n28922 , n19317 );
    and g18126 ( n19089 , n1741 , n7177 );
    not g18127 ( n6113 , n8054 );
    or g18128 ( n2396 , n2324 , n28241 );
    or g18129 ( n25046 , n13430 , n21967 );
    xnor g18130 ( n17324 , n22820 , n15642 );
    and g18131 ( n120 , n21555 , n2584 );
    nor g18132 ( n12252 , n1856 , n20390 );
    and g18133 ( n4464 , n22722 , n22945 );
    not g18134 ( n26259 , n664 );
    xnor g18135 ( n31792 , n22398 , n4997 );
    not g18136 ( n15928 , n5174 );
    not g18137 ( n13955 , n24697 );
    not g18138 ( n7341 , n19120 );
    not g18139 ( n26616 , n26139 );
    or g18140 ( n1390 , n139 , n22130 );
    and g18141 ( n12069 , n5461 , n24458 );
    not g18142 ( n12887 , n315 );
    not g18143 ( n14691 , n1012 );
    xnor g18144 ( n11527 , n13485 , n29604 );
    not g18145 ( n24388 , n8316 );
    and g18146 ( n29469 , n23662 , n12782 );
    xnor g18147 ( n27504 , n17227 , n27885 );
    or g18148 ( n23087 , n31019 , n18312 );
    buf g18149 ( n30238 , n19433 );
    xnor g18150 ( n22216 , n27245 , n11379 );
    not g18151 ( n31604 , n6136 );
    or g18152 ( n8010 , n10333 , n30202 );
    or g18153 ( n11748 , n6979 , n24376 );
    or g18154 ( n6771 , n20365 , n13733 );
    not g18155 ( n9983 , n27798 );
    not g18156 ( n28462 , n29466 );
    not g18157 ( n19939 , n18307 );
    or g18158 ( n28900 , n26665 , n9680 );
    xnor g18159 ( n16813 , n8574 , n6827 );
    and g18160 ( n10141 , n25899 , n1083 );
    or g18161 ( n20085 , n4417 , n9501 );
    not g18162 ( n24858 , n23683 );
    or g18163 ( n18433 , n14443 , n1823 );
    and g18164 ( n3862 , n1651 , n1620 );
    not g18165 ( n25016 , n30491 );
    nor g18166 ( n572 , n8005 , n30411 );
    or g18167 ( n23698 , n20220 , n15569 );
    not g18168 ( n16108 , n17617 );
    not g18169 ( n22615 , n8480 );
    or g18170 ( n6644 , n2098 , n20328 );
    nor g18171 ( n25686 , n24568 , n10152 );
    or g18172 ( n27819 , n27037 , n17246 );
    or g18173 ( n24927 , n31131 , n21405 );
    not g18174 ( n24382 , n22576 );
    not g18175 ( n4894 , n17025 );
    or g18176 ( n5798 , n20666 , n29491 );
    and g18177 ( n9365 , n15821 , n18270 );
    or g18178 ( n30725 , n272 , n18943 );
    xnor g18179 ( n6722 , n31450 , n6874 );
    or g18180 ( n6447 , n22625 , n18946 );
    xnor g18181 ( n21096 , n14180 , n24137 );
    not g18182 ( n14956 , n24697 );
    and g18183 ( n17610 , n96 , n25909 );
    not g18184 ( n27128 , n4997 );
    and g18185 ( n3247 , n10012 , n14725 );
    or g18186 ( n991 , n31203 , n28336 );
    and g18187 ( n31397 , n26760 , n26913 );
    not g18188 ( n25993 , n9300 );
    not g18189 ( n1207 , n18346 );
    nor g18190 ( n28420 , n29617 , n23249 );
    not g18191 ( n22777 , n21591 );
    xnor g18192 ( n6179 , n21925 , n16083 );
    xnor g18193 ( n9246 , n8501 , n22064 );
    buf g18194 ( n19524 , n6465 );
    and g18195 ( n4692 , n23149 , n17545 );
    not g18196 ( n198 , n4252 );
    nor g18197 ( n9381 , n9211 , n3787 );
    not g18198 ( n19142 , n138 );
    or g18199 ( n6215 , n18279 , n3773 );
    xnor g18200 ( n10961 , n19929 , n10608 );
    and g18201 ( n18428 , n26650 , n31941 );
    not g18202 ( n2246 , n20385 );
    xnor g18203 ( n8009 , n21884 , n2621 );
    nor g18204 ( n12878 , n2592 , n87 );
    not g18205 ( n26661 , n5800 );
    buf g18206 ( n3639 , n21591 );
    xnor g18207 ( n12245 , n3304 , n6915 );
    or g18208 ( n8892 , n15975 , n27820 );
    not g18209 ( n11640 , n9909 );
    and g18210 ( n26899 , n24556 , n253 );
    and g18211 ( n2166 , n31036 , n6728 );
    or g18212 ( n6458 , n14970 , n6083 );
    nor g18213 ( n2009 , n13840 , n16083 );
    not g18214 ( n20942 , n13382 );
    or g18215 ( n4871 , n30334 , n27016 );
    or g18216 ( n21254 , n28013 , n24489 );
    not g18217 ( n22792 , n23311 );
    xnor g18218 ( n6555 , n19472 , n12913 );
    not g18219 ( n29994 , n25227 );
    or g18220 ( n6933 , n3541 , n28133 );
    xnor g18221 ( n2337 , n29983 , n3619 );
    xnor g18222 ( n27113 , n8157 , n19743 );
    or g18223 ( n7850 , n18362 , n6211 );
    xnor g18224 ( n10977 , n14832 , n2911 );
    xnor g18225 ( n10322 , n15703 , n29968 );
    and g18226 ( n4018 , n24796 , n17939 );
    xnor g18227 ( n16098 , n4969 , n1360 );
    not g18228 ( n31175 , n13138 );
    nor g18229 ( n19748 , n3765 , n238 );
    not g18230 ( n1214 , n14835 );
    and g18231 ( n26972 , n26064 , n26892 );
    xnor g18232 ( n16708 , n28028 , n5083 );
    or g18233 ( n29652 , n4618 , n4571 );
    xnor g18234 ( n29031 , n1082 , n23992 );
    nor g18235 ( n10813 , n22451 , n3973 );
    or g18236 ( n15314 , n32033 , n28513 );
    not g18237 ( n24141 , n3420 );
    or g18238 ( n19219 , n19615 , n5906 );
    not g18239 ( n31855 , n25755 );
    and g18240 ( n25060 , n10715 , n5074 );
    xnor g18241 ( n14545 , n2188 , n26746 );
    not g18242 ( n27409 , n9689 );
    or g18243 ( n21837 , n6837 , n27697 );
    or g18244 ( n15241 , n8662 , n21777 );
    or g18245 ( n31827 , n9871 , n16068 );
    not g18246 ( n1117 , n27213 );
    or g18247 ( n31692 , n25132 , n20605 );
    or g18248 ( n29634 , n17910 , n11248 );
    or g18249 ( n27727 , n15588 , n16075 );
    xnor g18250 ( n23886 , n2376 , n30084 );
    not g18251 ( n30383 , n11344 );
    not g18252 ( n28384 , n28452 );
    not g18253 ( n30268 , n11372 );
    xnor g18254 ( n11355 , n15781 , n20125 );
    nor g18255 ( n14315 , n4916 , n3949 );
    not g18256 ( n13122 , n18035 );
    or g18257 ( n26781 , n26983 , n22753 );
    or g18258 ( n9614 , n16237 , n12551 );
    not g18259 ( n27109 , n408 );
    and g18260 ( n11377 , n27725 , n28529 );
    not g18261 ( n15447 , n21036 );
    or g18262 ( n10993 , n201 , n5577 );
    or g18263 ( n30774 , n27273 , n23404 );
    or g18264 ( n22547 , n24121 , n19441 );
    not g18265 ( n10467 , n5125 );
    not g18266 ( n27215 , n9418 );
    xnor g18267 ( n11279 , n3254 , n9016 );
    or g18268 ( n24200 , n6466 , n5791 );
    not g18269 ( n14836 , n26882 );
    not g18270 ( n31549 , n11450 );
    not g18271 ( n29187 , n3157 );
    xnor g18272 ( n4652 , n25585 , n18165 );
    xnor g18273 ( n3511 , n27896 , n11610 );
    xnor g18274 ( n29655 , n16186 , n20603 );
    buf g18275 ( n24008 , n17141 );
    not g18276 ( n22069 , n27646 );
    not g18277 ( n30490 , n19642 );
    xnor g18278 ( n25693 , n22907 , n21104 );
    nor g18279 ( n9623 , n11598 , n22022 );
    nor g18280 ( n12749 , n16873 , n6084 );
    not g18281 ( n4915 , n10599 );
    xor g18282 ( n25557 , n17748 , n3985 );
    xnor g18283 ( n11702 , n2939 , n12514 );
    and g18284 ( n8142 , n29675 , n20547 );
    or g18285 ( n9562 , n11575 , n25655 );
    not g18286 ( n25422 , n17457 );
    or g18287 ( n12152 , n20027 , n14862 );
    xnor g18288 ( n9060 , n18036 , n16376 );
    or g18289 ( n28826 , n22233 , n25300 );
    or g18290 ( n9848 , n22260 , n8250 );
    not g18291 ( n12439 , n19317 );
    not g18292 ( n24977 , n7349 );
    xnor g18293 ( n30894 , n21740 , n17872 );
    xnor g18294 ( n6550 , n16126 , n17885 );
    xnor g18295 ( n17783 , n29957 , n5914 );
    or g18296 ( n2682 , n15731 , n20068 );
    not g18297 ( n14014 , n11642 );
    and g18298 ( n29477 , n11878 , n14365 );
    xnor g18299 ( n22525 , n10023 , n16058 );
    xnor g18300 ( n6380 , n27515 , n13150 );
    nor g18301 ( n6515 , n6251 , n6881 );
    xnor g18302 ( n3859 , n23898 , n4790 );
    and g18303 ( n15291 , n19415 , n29175 );
    and g18304 ( n27659 , n31630 , n31574 );
    xnor g18305 ( n1455 , n14015 , n6751 );
    or g18306 ( n20816 , n3265 , n26998 );
    xnor g18307 ( n14958 , n16258 , n21381 );
    xnor g18308 ( n2191 , n17068 , n11218 );
    or g18309 ( n18894 , n21597 , n12428 );
    xnor g18310 ( n22909 , n12538 , n18473 );
    nor g18311 ( n19535 , n8809 , n23337 );
    nor g18312 ( n22824 , n30158 , n25242 );
    or g18313 ( n15707 , n28180 , n11517 );
    xnor g18314 ( n10193 , n17962 , n3096 );
    nor g18315 ( n23354 , n19561 , n27221 );
    xnor g18316 ( n9531 , n21236 , n31654 );
    and g18317 ( n27307 , n13174 , n5338 );
    or g18318 ( n29104 , n4501 , n10046 );
    xnor g18319 ( n30805 , n23191 , n20939 );
    nor g18320 ( n26234 , n18253 , n13281 );
    xnor g18321 ( n18438 , n10501 , n9502 );
    xnor g18322 ( n29662 , n15120 , n12798 );
    not g18323 ( n31873 , n22204 );
    and g18324 ( n10138 , n13177 , n30967 );
    xnor g18325 ( n961 , n2366 , n27792 );
    and g18326 ( n1970 , n4834 , n3904 );
    and g18327 ( n1329 , n11985 , n23391 );
    and g18328 ( n28423 , n11079 , n24491 );
    xnor g18329 ( n21531 , n14872 , n29668 );
    or g18330 ( n16253 , n3032 , n21240 );
    not g18331 ( n3939 , n13201 );
    and g18332 ( n15426 , n8226 , n500 );
    xnor g18333 ( n276 , n19084 , n214 );
    or g18334 ( n13584 , n11197 , n27184 );
    xnor g18335 ( n9580 , n2267 , n21392 );
    and g18336 ( n9221 , n1324 , n5160 );
    not g18337 ( n1097 , n30557 );
    or g18338 ( n29868 , n20184 , n4289 );
    not g18339 ( n12 , n16203 );
    not g18340 ( n21514 , n27251 );
    nor g18341 ( n11665 , n9795 , n11382 );
    xnor g18342 ( n20026 , n18902 , n117 );
    not g18343 ( n25056 , n8269 );
    not g18344 ( n29779 , n22902 );
    nor g18345 ( n1169 , n3269 , n7103 );
    xnor g18346 ( n31007 , n4078 , n20811 );
    and g18347 ( n29263 , n18594 , n2341 );
    or g18348 ( n9171 , n6277 , n20645 );
    buf g18349 ( n346 , n8330 );
    or g18350 ( n25451 , n31791 , n20268 );
    xnor g18351 ( n20805 , n11851 , n18389 );
    and g18352 ( n22437 , n1832 , n24548 );
    or g18353 ( n8373 , n22858 , n25980 );
    and g18354 ( n8141 , n29342 , n27899 );
    or g18355 ( n21985 , n26490 , n28027 );
    not g18356 ( n28678 , n29706 );
    or g18357 ( n7297 , n27594 , n3589 );
    xnor g18358 ( n18393 , n20216 , n11155 );
    not g18359 ( n580 , n18381 );
    xnor g18360 ( n19712 , n561 , n29132 );
    xnor g18361 ( n19443 , n25528 , n5046 );
    or g18362 ( n21713 , n5806 , n2288 );
    or g18363 ( n5647 , n19592 , n24852 );
    and g18364 ( n1497 , n24971 , n28120 );
    or g18365 ( n12236 , n23814 , n27795 );
    xnor g18366 ( n13440 , n11218 , n2447 );
    xnor g18367 ( n5922 , n841 , n22726 );
    not g18368 ( n5058 , n29326 );
    or g18369 ( n25922 , n20993 , n20628 );
    or g18370 ( n14529 , n7412 , n7751 );
    or g18371 ( n10303 , n9691 , n32021 );
    and g18372 ( n8911 , n11451 , n10885 );
    and g18373 ( n22219 , n1777 , n26773 );
    xnor g18374 ( n13835 , n12920 , n8713 );
    not g18375 ( n25720 , n26494 );
    not g18376 ( n221 , n21410 );
    not g18377 ( n302 , n26894 );
    not g18378 ( n23676 , n27829 );
    and g18379 ( n7382 , n17516 , n29257 );
    and g18380 ( n24979 , n18050 , n1399 );
    or g18381 ( n1805 , n13938 , n27875 );
    or g18382 ( n29220 , n23743 , n7956 );
    nor g18383 ( n9045 , n3131 , n20881 );
    not g18384 ( n28578 , n23788 );
    or g18385 ( n30592 , n25325 , n20678 );
    or g18386 ( n1838 , n23232 , n16414 );
    nor g18387 ( n15843 , n13865 , n13267 );
    xnor g18388 ( n18670 , n5389 , n17172 );
    xnor g18389 ( n14769 , n31271 , n19282 );
    not g18390 ( n28020 , n12845 );
    not g18391 ( n7497 , n29870 );
    or g18392 ( n30078 , n18938 , n8444 );
    or g18393 ( n4100 , n7692 , n4848 );
    and g18394 ( n11885 , n27001 , n5908 );
    or g18395 ( n29713 , n3403 , n13089 );
    nor g18396 ( n27331 , n30326 , n28736 );
    not g18397 ( n2243 , n19915 );
    or g18398 ( n13258 , n1610 , n8779 );
    not g18399 ( n3938 , n28787 );
    and g18400 ( n20450 , n3742 , n9392 );
    or g18401 ( n5051 , n19908 , n22409 );
    and g18402 ( n14382 , n26086 , n24551 );
    and g18403 ( n12881 , n19606 , n9649 );
    or g18404 ( n6684 , n25339 , n19822 );
    or g18405 ( n20263 , n11771 , n1696 );
    xnor g18406 ( n27370 , n18100 , n19187 );
    xnor g18407 ( n14257 , n16885 , n5310 );
    xnor g18408 ( n2486 , n10708 , n172 );
    or g18409 ( n9997 , n24358 , n17298 );
    xnor g18410 ( n14851 , n20236 , n17843 );
    or g18411 ( n5795 , n8835 , n2859 );
    xnor g18412 ( n16110 , n21235 , n27354 );
    or g18413 ( n11769 , n25174 , n3069 );
    and g18414 ( n31123 , n24181 , n2331 );
    xnor g18415 ( n21707 , n24071 , n7063 );
    or g18416 ( n5877 , n17109 , n25728 );
    and g18417 ( n11241 , n15090 , n15427 );
    not g18418 ( n5518 , n7879 );
    xnor g18419 ( n24822 , n3993 , n12105 );
    nor g18420 ( n20273 , n17343 , n13950 );
    xnor g18421 ( n19622 , n23237 , n29050 );
    not g18422 ( n5749 , n21156 );
    not g18423 ( n8538 , n24358 );
    or g18424 ( n4123 , n27094 , n23224 );
    and g18425 ( n22834 , n15712 , n7166 );
    xnor g18426 ( n2764 , n28237 , n29878 );
    xnor g18427 ( n15870 , n11205 , n29090 );
    or g18428 ( n333 , n22517 , n8671 );
    or g18429 ( n1409 , n13454 , n8014 );
    or g18430 ( n21069 , n7785 , n20606 );
    or g18431 ( n26398 , n6285 , n4955 );
    or g18432 ( n4598 , n15853 , n3159 );
    xor g18433 ( n16260 , n5869 , n6940 );
    xnor g18434 ( n31633 , n6651 , n2150 );
    nor g18435 ( n27182 , n16836 , n17684 );
    xor g18436 ( n4777 , n1877 , n3341 );
    and g18437 ( n13824 , n10531 , n26431 );
    not g18438 ( n21417 , n13676 );
    or g18439 ( n27642 , n5150 , n5873 );
    xnor g18440 ( n17550 , n30884 , n1893 );
    xnor g18441 ( n17501 , n12437 , n31338 );
    nor g18442 ( n4294 , n20274 , n5045 );
    xnor g18443 ( n9428 , n5774 , n241 );
    nor g18444 ( n28991 , n21653 , n13425 );
    or g18445 ( n27387 , n11658 , n21995 );
    not g18446 ( n25393 , n9531 );
    xnor g18447 ( n25333 , n27918 , n16493 );
    xnor g18448 ( n9776 , n25128 , n18015 );
    not g18449 ( n19472 , n15391 );
    xnor g18450 ( n18298 , n3166 , n18394 );
    and g18451 ( n1000 , n8334 , n3275 );
    not g18452 ( n10105 , n21603 );
    not g18453 ( n14510 , n27019 );
    xnor g18454 ( n27615 , n19899 , n1483 );
    not g18455 ( n28666 , n22570 );
    xnor g18456 ( n12020 , n14495 , n27439 );
    or g18457 ( n24373 , n3303 , n4610 );
    not g18458 ( n7820 , n21480 );
    or g18459 ( n7916 , n19098 , n15247 );
    not g18460 ( n6302 , n30167 );
    and g18461 ( n13474 , n23445 , n5505 );
    not g18462 ( n8580 , n13973 );
    xnor g18463 ( n24047 , n23352 , n25768 );
    or g18464 ( n18144 , n14391 , n20473 );
    and g18465 ( n29155 , n19286 , n2478 );
    xnor g18466 ( n22167 , n30978 , n16071 );
    xnor g18467 ( n20031 , n17303 , n27298 );
    not g18468 ( n3710 , n3829 );
    nor g18469 ( n15681 , n13975 , n30853 );
    xnor g18470 ( n2316 , n31317 , n14825 );
    or g18471 ( n15481 , n4847 , n25643 );
    xnor g18472 ( n22223 , n9310 , n4924 );
    not g18473 ( n1718 , n31616 );
    nor g18474 ( n16764 , n22845 , n18507 );
    xnor g18475 ( n24767 , n26274 , n28965 );
    not g18476 ( n17032 , n26598 );
    not g18477 ( n16956 , n11756 );
    xnor g18478 ( n27090 , n26913 , n26760 );
    nor g18479 ( n27372 , n2825 , n1604 );
    xor g18480 ( n16010 , n24193 , n14386 );
    or g18481 ( n1514 , n25272 , n21166 );
    xnor g18482 ( n25726 , n7360 , n1123 );
    xnor g18483 ( n5377 , n5186 , n26606 );
    and g18484 ( n25647 , n20748 , n30287 );
    or g18485 ( n10829 , n12373 , n6453 );
    not g18486 ( n10097 , n1120 );
    or g18487 ( n12909 , n16318 , n31841 );
    and g18488 ( n3632 , n9488 , n8804 );
    not g18489 ( n7746 , n12279 );
    not g18490 ( n29637 , n6881 );
    or g18491 ( n8069 , n7303 , n7889 );
    or g18492 ( n21699 , n25757 , n7999 );
    not g18493 ( n21932 , n19434 );
    or g18494 ( n25232 , n1746 , n9395 );
    and g18495 ( n17738 , n27518 , n31872 );
    not g18496 ( n18286 , n8579 );
    not g18497 ( n12953 , n25259 );
    xnor g18498 ( n14016 , n17581 , n10932 );
    xor g18499 ( n2542 , n16898 , n17417 );
    or g18500 ( n57 , n9572 , n9057 );
    or g18501 ( n9136 , n10576 , n22486 );
    xnor g18502 ( n4182 , n24650 , n28139 );
    and g18503 ( n19293 , n26442 , n23211 );
    not g18504 ( n20146 , n13467 );
    xnor g18505 ( n3040 , n13690 , n22349 );
    and g18506 ( n8463 , n10341 , n1778 );
    xnor g18507 ( n28587 , n22759 , n18534 );
    or g18508 ( n30050 , n10580 , n27437 );
    or g18509 ( n27337 , n23971 , n8199 );
    and g18510 ( n14340 , n1900 , n9289 );
    or g18511 ( n19851 , n1854 , n15308 );
    not g18512 ( n5528 , n10871 );
    xnor g18513 ( n17613 , n15830 , n3795 );
    xnor g18514 ( n16227 , n1831 , n6534 );
    not g18515 ( n20755 , n31563 );
    nor g18516 ( n29164 , n18612 , n2473 );
    or g18517 ( n20925 , n12965 , n12191 );
    not g18518 ( n14196 , n8602 );
    xnor g18519 ( n27396 , n1300 , n12287 );
    xnor g18520 ( n29053 , n21128 , n7864 );
    not g18521 ( n7662 , n17974 );
    xnor g18522 ( n13338 , n12107 , n31348 );
    xnor g18523 ( n31702 , n569 , n21945 );
    xnor g18524 ( n14519 , n13970 , n1429 );
    nor g18525 ( n18891 , n21507 , n26047 );
    xnor g18526 ( n28326 , n2817 , n10884 );
    or g18527 ( n1392 , n15242 , n21281 );
    or g18528 ( n19555 , n4213 , n20171 );
    nor g18529 ( n23494 , n26863 , n9402 );
    xnor g18530 ( n19212 , n4002 , n4124 );
    or g18531 ( n28710 , n25684 , n6520 );
    not g18532 ( n29218 , n2020 );
    or g18533 ( n17935 , n31889 , n28470 );
    not g18534 ( n29466 , n9005 );
    not g18535 ( n30000 , n4571 );
    xnor g18536 ( n17304 , n7314 , n8321 );
    buf g18537 ( n10713 , n30394 );
    not g18538 ( n29991 , n3906 );
    nor g18539 ( n21599 , n23052 , n579 );
    or g18540 ( n30662 , n19741 , n22789 );
    or g18541 ( n25540 , n9613 , n10084 );
    or g18542 ( n7275 , n4091 , n3675 );
    and g18543 ( n1055 , n25604 , n12679 );
    xnor g18544 ( n17461 , n20632 , n20759 );
    or g18545 ( n1547 , n27695 , n4789 );
    and g18546 ( n2780 , n2613 , n15993 );
    or g18547 ( n15541 , n24880 , n6621 );
    or g18548 ( n20699 , n8005 , n777 );
    not g18549 ( n18281 , n14298 );
    xnor g18550 ( n89 , n19231 , n17851 );
    xnor g18551 ( n27080 , n11993 , n9691 );
    not g18552 ( n8282 , n13022 );
    or g18553 ( n7953 , n28611 , n12893 );
    or g18554 ( n2729 , n2997 , n14821 );
    xnor g18555 ( n11653 , n2419 , n4209 );
    or g18556 ( n12667 , n3038 , n23356 );
    not g18557 ( n21472 , n10200 );
    and g18558 ( n17669 , n3429 , n18303 );
    or g18559 ( n25039 , n17063 , n1807 );
    not g18560 ( n4778 , n18418 );
    and g18561 ( n21042 , n5666 , n24140 );
    xor g18562 ( n22235 , n14472 , n25924 );
    and g18563 ( n4036 , n3212 , n31678 );
    not g18564 ( n6014 , n4814 );
    and g18565 ( n1842 , n29411 , n28734 );
    not g18566 ( n7880 , n8654 );
    and g18567 ( n14182 , n13159 , n10405 );
    not g18568 ( n5814 , n11610 );
    and g18569 ( n4329 , n8193 , n915 );
    and g18570 ( n20899 , n26402 , n6468 );
    or g18571 ( n21590 , n9836 , n2042 );
    xnor g18572 ( n11227 , n7042 , n25255 );
    not g18573 ( n10700 , n5982 );
    not g18574 ( n16851 , n5848 );
    nor g18575 ( n9165 , n6626 , n14537 );
    not g18576 ( n8403 , n13700 );
    not g18577 ( n1316 , n22113 );
    or g18578 ( n26900 , n31121 , n7597 );
    nor g18579 ( n1976 , n12428 , n4480 );
    or g18580 ( n5311 , n24680 , n30333 );
    buf g18581 ( n10196 , n20480 );
    or g18582 ( n4178 , n12665 , n21499 );
    or g18583 ( n915 , n26 , n13249 );
    xnor g18584 ( n3590 , n14937 , n25674 );
    xnor g18585 ( n26242 , n13800 , n2629 );
    xnor g18586 ( n25049 , n1326 , n15260 );
    nor g18587 ( n24199 , n26871 , n9104 );
    or g18588 ( n19806 , n19942 , n16362 );
    xnor g18589 ( n22194 , n6969 , n22902 );
    and g18590 ( n20399 , n28710 , n14113 );
    xnor g18591 ( n4958 , n17433 , n22826 );
    and g18592 ( n10886 , n22468 , n9312 );
    not g18593 ( n3033 , n7762 );
    xnor g18594 ( n20703 , n3752 , n6483 );
    not g18595 ( n30429 , n24164 );
    xnor g18596 ( n21076 , n13704 , n23400 );
    not g18597 ( n31491 , n7928 );
    not g18598 ( n672 , n5792 );
    xnor g18599 ( n14571 , n7415 , n7464 );
    and g18600 ( n30618 , n27672 , n24212 );
    or g18601 ( n4413 , n19096 , n16757 );
    not g18602 ( n3867 , n5690 );
    nor g18603 ( n29370 , n3762 , n24468 );
    not g18604 ( n6970 , n1742 );
    xnor g18605 ( n25157 , n20033 , n26218 );
    or g18606 ( n8105 , n14767 , n14281 );
    nor g18607 ( n16664 , n13734 , n4813 );
    nor g18608 ( n21542 , n2883 , n16340 );
    xnor g18609 ( n1712 , n13448 , n8873 );
    not g18610 ( n6494 , n26198 );
    not g18611 ( n5126 , n1057 );
    xnor g18612 ( n29452 , n3100 , n29542 );
    or g18613 ( n28418 , n24768 , n24372 );
    nor g18614 ( n9225 , n4554 , n31889 );
    and g18615 ( n15381 , n2122 , n11856 );
    xnor g18616 ( n4665 , n11723 , n7648 );
    or g18617 ( n14032 , n20821 , n15290 );
    xnor g18618 ( n22464 , n16347 , n12627 );
    xnor g18619 ( n25248 , n26982 , n4069 );
    xnor g18620 ( n13029 , n6956 , n21346 );
    xnor g18621 ( n802 , n28721 , n16171 );
    nor g18622 ( n916 , n22595 , n31393 );
    not g18623 ( n1894 , n18350 );
    nor g18624 ( n11212 , n20156 , n23138 );
    nor g18625 ( n22055 , n30572 , n13989 );
    not g18626 ( n51 , n23483 );
    or g18627 ( n16388 , n4197 , n11268 );
    and g18628 ( n4241 , n26013 , n27984 );
    nor g18629 ( n7146 , n15530 , n12488 );
    and g18630 ( n21955 , n5763 , n3960 );
    xnor g18631 ( n23094 , n24821 , n29620 );
    not g18632 ( n2135 , n6858 );
    and g18633 ( n19954 , n25205 , n10650 );
    not g18634 ( n28998 , n6974 );
    not g18635 ( n30784 , n9398 );
    and g18636 ( n19729 , n7590 , n8548 );
    xnor g18637 ( n13834 , n13036 , n30941 );
    xnor g18638 ( n17293 , n23274 , n11380 );
    xnor g18639 ( n8200 , n24967 , n23970 );
    nor g18640 ( n23134 , n25291 , n15638 );
    not g18641 ( n27783 , n23348 );
    xnor g18642 ( n31686 , n2025 , n16191 );
    or g18643 ( n21958 , n221 , n15144 );
    and g18644 ( n29648 , n25157 , n10196 );
    nor g18645 ( n27850 , n1178 , n22154 );
    not g18646 ( n17542 , n24355 );
    or g18647 ( n26630 , n26664 , n31239 );
    not g18648 ( n7843 , n17306 );
    not g18649 ( n11605 , n24613 );
    xnor g18650 ( n15846 , n27327 , n21276 );
    not g18651 ( n30785 , n10081 );
    not g18652 ( n25682 , n22307 );
    or g18653 ( n20733 , n147 , n3950 );
    or g18654 ( n17770 , n9250 , n4581 );
    or g18655 ( n22769 , n23760 , n5777 );
    not g18656 ( n5078 , n23561 );
    not g18657 ( n9812 , n3661 );
    xnor g18658 ( n11906 , n6050 , n10522 );
    xnor g18659 ( n10774 , n6863 , n31924 );
    not g18660 ( n26611 , n2648 );
    or g18661 ( n21905 , n5939 , n17976 );
    and g18662 ( n21877 , n22926 , n26394 );
    or g18663 ( n16016 , n20329 , n28596 );
    xnor g18664 ( n17473 , n20576 , n10242 );
    nor g18665 ( n24228 , n17917 , n25167 );
    xnor g18666 ( n26849 , n1098 , n20756 );
    not g18667 ( n29065 , n4754 );
    xnor g18668 ( n26573 , n30099 , n1593 );
    xnor g18669 ( n7163 , n25294 , n15863 );
    and g18670 ( n19181 , n17340 , n25080 );
    or g18671 ( n6799 , n8013 , n6126 );
    and g18672 ( n15488 , n18915 , n8705 );
    not g18673 ( n30121 , n27738 );
    and g18674 ( n8694 , n18083 , n14355 );
    nor g18675 ( n11953 , n13800 , n12524 );
    nor g18676 ( n15014 , n3163 , n1036 );
    not g18677 ( n8572 , n24520 );
    nor g18678 ( n7367 , n23419 , n20046 );
    not g18679 ( n23644 , n3564 );
    nor g18680 ( n11802 , n28081 , n3509 );
    xnor g18681 ( n23068 , n22549 , n17499 );
    xnor g18682 ( n7047 , n611 , n30279 );
    not g18683 ( n15678 , n5898 );
    not g18684 ( n15310 , n21953 );
    and g18685 ( n2857 , n30263 , n19583 );
    xnor g18686 ( n6160 , n28267 , n6651 );
    not g18687 ( n5838 , n23330 );
    xnor g18688 ( n22956 , n10688 , n10776 );
    not g18689 ( n14731 , n20962 );
    not g18690 ( n7172 , n3793 );
    xnor g18691 ( n3030 , n7858 , n9244 );
    xnor g18692 ( n5449 , n12639 , n3480 );
    xnor g18693 ( n21470 , n26917 , n20042 );
    not g18694 ( n25261 , n24795 );
    not g18695 ( n2296 , n6650 );
    or g18696 ( n30637 , n27723 , n15462 );
    xnor g18697 ( n26656 , n8577 , n22867 );
    and g18698 ( n2036 , n24475 , n8652 );
    or g18699 ( n25998 , n31544 , n24899 );
    not g18700 ( n12212 , n19143 );
    or g18701 ( n29088 , n6048 , n20340 );
    and g18702 ( n29169 , n13388 , n31202 );
    or g18703 ( n11113 , n21461 , n10720 );
    nor g18704 ( n12274 , n23648 , n3567 );
    not g18705 ( n30893 , n21373 );
    xnor g18706 ( n31534 , n28037 , n10925 );
    not g18707 ( n30006 , n7729 );
    not g18708 ( n14643 , n16019 );
    xnor g18709 ( n27833 , n15961 , n26796 );
    or g18710 ( n5971 , n6256 , n16277 );
    or g18711 ( n25381 , n29679 , n22407 );
    nor g18712 ( n8149 , n3677 , n4507 );
    and g18713 ( n1548 , n2197 , n29713 );
    not g18714 ( n6381 , n6445 );
    or g18715 ( n12483 , n28401 , n30137 );
    not g18716 ( n31435 , n10393 );
    nor g18717 ( n17206 , n22917 , n785 );
    xnor g18718 ( n16055 , n30343 , n3163 );
    or g18719 ( n7954 , n24647 , n15808 );
    or g18720 ( n25185 , n20154 , n8120 );
    not g18721 ( n5839 , n22617 );
    not g18722 ( n10952 , n31773 );
    or g18723 ( n19329 , n10482 , n9117 );
    xnor g18724 ( n27973 , n26219 , n29938 );
    not g18725 ( n9920 , n21257 );
    or g18726 ( n22784 , n7669 , n23461 );
    nor g18727 ( n25505 , n19231 , n4358 );
    not g18728 ( n12054 , n29525 );
    xnor g18729 ( n30800 , n24899 , n14713 );
    and g18730 ( n29606 , n18604 , n20116 );
    xnor g18731 ( n2392 , n18828 , n6510 );
    not g18732 ( n12123 , n22576 );
    and g18733 ( n2952 , n17608 , n25965 );
    buf g18734 ( n31595 , n7796 );
    or g18735 ( n29277 , n8014 , n13402 );
    or g18736 ( n23429 , n13255 , n26589 );
    not g18737 ( n9208 , n12060 );
    xnor g18738 ( n22721 , n165 , n19869 );
    and g18739 ( n19497 , n18670 , n14276 );
    and g18740 ( n6002 , n27998 , n9968 );
    not g18741 ( n30642 , n16586 );
    nor g18742 ( n5784 , n6888 , n21084 );
    nor g18743 ( n19918 , n6191 , n22802 );
    not g18744 ( n5222 , n24824 );
    or g18745 ( n17383 , n21759 , n12537 );
    xnor g18746 ( n28719 , n22114 , n8852 );
    not g18747 ( n31885 , n28951 );
    or g18748 ( n10189 , n2401 , n21505 );
    xnor g18749 ( n29070 , n20542 , n14189 );
    and g18750 ( n5671 , n31444 , n29067 );
    xnor g18751 ( n17127 , n4426 , n4701 );
    not g18752 ( n29664 , n16145 );
    or g18753 ( n21737 , n21272 , n17342 );
    not g18754 ( n19343 , n19943 );
    xnor g18755 ( n5060 , n9869 , n18252 );
    or g18756 ( n8148 , n4725 , n8459 );
    xnor g18757 ( n19206 , n9914 , n18518 );
    xnor g18758 ( n25678 , n30025 , n12777 );
    not g18759 ( n21911 , n18255 );
    or g18760 ( n12834 , n17815 , n25401 );
    not g18761 ( n20774 , n7491 );
    or g18762 ( n28760 , n8831 , n10381 );
    xor g18763 ( n3668 , n22982 , n19193 );
    and g18764 ( n22323 , n8154 , n6113 );
    not g18765 ( n5688 , n6535 );
    not g18766 ( n6026 , n5628 );
    nor g18767 ( n17134 , n13175 , n11147 );
    xnor g18768 ( n17986 , n16581 , n24667 );
    nor g18769 ( n12361 , n18438 , n21893 );
    and g18770 ( n13357 , n11475 , n25186 );
    xnor g18771 ( n9785 , n10500 , n10407 );
    and g18772 ( n23371 , n1726 , n28352 );
    not g18773 ( n1755 , n12131 );
    and g18774 ( n16116 , n2976 , n31249 );
    and g18775 ( n10323 , n13227 , n1547 );
    xnor g18776 ( n24311 , n25062 , n3439 );
    or g18777 ( n12010 , n2798 , n31635 );
    not g18778 ( n3558 , n16233 );
    and g18779 ( n30965 , n13586 , n27938 );
    and g18780 ( n16517 , n8730 , n6563 );
    not g18781 ( n12444 , n7891 );
    not g18782 ( n21595 , n7057 );
    not g18783 ( n7378 , n24335 );
    or g18784 ( n31814 , n23016 , n6724 );
    not g18785 ( n10435 , n14925 );
    xnor g18786 ( n22742 , n21960 , n23047 );
    not g18787 ( n30466 , n31761 );
    and g18788 ( n24505 , n15018 , n16451 );
    not g18789 ( n28549 , n22626 );
    or g18790 ( n801 , n16294 , n12473 );
    or g18791 ( n3044 , n11171 , n16248 );
    not g18792 ( n10222 , n29093 );
    xnor g18793 ( n28975 , n31901 , n16774 );
    not g18794 ( n16872 , n27872 );
    not g18795 ( n11412 , n27615 );
    not g18796 ( n25353 , n17890 );
    not g18797 ( n6985 , n16760 );
    and g18798 ( n25575 , n2807 , n19527 );
    and g18799 ( n705 , n22653 , n3712 );
    and g18800 ( n8476 , n26611 , n3637 );
    not g18801 ( n7715 , n30871 );
    xnor g18802 ( n18908 , n12065 , n24415 );
    xnor g18803 ( n17082 , n6750 , n21180 );
    nor g18804 ( n10668 , n31856 , n23823 );
    xnor g18805 ( n3571 , n13145 , n29437 );
    or g18806 ( n18665 , n24939 , n26395 );
    xnor g18807 ( n4300 , n3473 , n26418 );
    or g18808 ( n25294 , n28505 , n23467 );
    xnor g18809 ( n5898 , n16899 , n7101 );
    xnor g18810 ( n26764 , n30012 , n29981 );
    and g18811 ( n16160 , n21121 , n22764 );
    or g18812 ( n27739 , n9842 , n25237 );
    and g18813 ( n14462 , n26039 , n14265 );
    xnor g18814 ( n919 , n23428 , n9891 );
    or g18815 ( n21975 , n962 , n20126 );
    buf g18816 ( n6046 , n26676 );
    or g18817 ( n1456 , n26797 , n9106 );
    xor g18818 ( n12384 , n24796 , n18701 );
    xnor g18819 ( n5170 , n6629 , n26267 );
    xnor g18820 ( n20591 , n832 , n20227 );
    nor g18821 ( n13144 , n31404 , n8705 );
    and g18822 ( n26562 , n20668 , n28038 );
    xnor g18823 ( n718 , n25748 , n5637 );
    nor g18824 ( n8618 , n15166 , n17334 );
    xnor g18825 ( n13850 , n16829 , n3800 );
    not g18826 ( n5675 , n21174 );
    and g18827 ( n15093 , n20054 , n6588 );
    xnor g18828 ( n5721 , n29577 , n27981 );
    xnor g18829 ( n31647 , n1094 , n21469 );
    or g18830 ( n3309 , n25101 , n356 );
    nor g18831 ( n14381 , n24884 , n10597 );
    nor g18832 ( n23324 , n14872 , n8255 );
    not g18833 ( n30874 , n22369 );
    xnor g18834 ( n25234 , n25297 , n11253 );
    and g18835 ( n7807 , n30382 , n20670 );
    xnor g18836 ( n11269 , n2143 , n11770 );
    xnor g18837 ( n31736 , n24813 , n6106 );
    and g18838 ( n24486 , n9849 , n31801 );
    not g18839 ( n2936 , n13657 );
    and g18840 ( n23432 , n2456 , n13027 );
    not g18841 ( n4859 , n17261 );
    not g18842 ( n18912 , n18442 );
    and g18843 ( n17153 , n27809 , n25908 );
    and g18844 ( n30151 , n31766 , n22704 );
    not g18845 ( n13535 , n19615 );
    and g18846 ( n6892 , n11398 , n30197 );
    or g18847 ( n24541 , n31234 , n18934 );
    not g18848 ( n27238 , n29984 );
    not g18849 ( n20335 , n29777 );
    nor g18850 ( n6218 , n5202 , n26193 );
    not g18851 ( n31026 , n13744 );
    and g18852 ( n13868 , n8819 , n8308 );
    not g18853 ( n14936 , n19615 );
    not g18854 ( n7763 , n25491 );
    nor g18855 ( n27677 , n5271 , n22248 );
    xnor g18856 ( n30444 , n12367 , n29909 );
    or g18857 ( n8254 , n8873 , n28501 );
    not g18858 ( n12011 , n18775 );
    xnor g18859 ( n5442 , n27078 , n7657 );
    or g18860 ( n46 , n19121 , n21927 );
    or g18861 ( n30609 , n4164 , n14349 );
    and g18862 ( n9106 , n693 , n1925 );
    not g18863 ( n28616 , n42 );
    and g18864 ( n5743 , n14158 , n18777 );
    or g18865 ( n9839 , n17898 , n30997 );
    xnor g18866 ( n1348 , n28421 , n15370 );
    not g18867 ( n24143 , n6720 );
    or g18868 ( n29758 , n5403 , n19815 );
    or g18869 ( n18573 , n8914 , n21295 );
    nor g18870 ( n17868 , n18808 , n16292 );
    nor g18871 ( n14905 , n31970 , n9053 );
    not g18872 ( n1797 , n14943 );
    not g18873 ( n17131 , n9208 );
    xnor g18874 ( n16938 , n16806 , n27690 );
    or g18875 ( n12776 , n3632 , n10412 );
    not g18876 ( n19564 , n8195 );
    not g18877 ( n21399 , n26746 );
    and g18878 ( n15854 , n11559 , n30175 );
    xnor g18879 ( n4849 , n24614 , n20031 );
    or g18880 ( n13306 , n30245 , n1600 );
    xnor g18881 ( n23336 , n4323 , n5379 );
    or g18882 ( n4938 , n21957 , n15597 );
    or g18883 ( n6444 , n19598 , n16398 );
    not g18884 ( n4454 , n2236 );
    buf g18885 ( n10955 , n10082 );
    not g18886 ( n1093 , n5818 );
    xnor g18887 ( n4833 , n20013 , n8901 );
    not g18888 ( n12609 , n23776 );
    or g18889 ( n6531 , n13302 , n5264 );
    not g18890 ( n17474 , n12630 );
    and g18891 ( n13482 , n11639 , n31679 );
    nor g18892 ( n12487 , n31727 , n7354 );
    xor g18893 ( n23032 , n6104 , n29173 );
    not g18894 ( n23083 , n31337 );
    or g18895 ( n30653 , n4109 , n16668 );
    not g18896 ( n12246 , n20514 );
    nor g18897 ( n24034 , n2934 , n25063 );
    or g18898 ( n10783 , n2486 , n8845 );
    nor g18899 ( n21457 , n25585 , n18165 );
    xnor g18900 ( n29660 , n18585 , n30706 );
    xor g18901 ( n25144 , n7885 , n18376 );
    and g18902 ( n7686 , n20073 , n18982 );
    nor g18903 ( n22271 , n16725 , n26325 );
    xnor g18904 ( n22454 , n14281 , n6971 );
    nor g18905 ( n24024 , n21736 , n1278 );
    and g18906 ( n25779 , n318 , n14489 );
    and g18907 ( n17154 , n19217 , n21136 );
    not g18908 ( n2981 , n27591 );
    or g18909 ( n611 , n1391 , n8765 );
    or g18910 ( n28493 , n12803 , n29368 );
    or g18911 ( n27257 , n17380 , n416 );
    not g18912 ( n9037 , n15076 );
    not g18913 ( n30313 , n23474 );
    not g18914 ( n3490 , n16986 );
    nor g18915 ( n26453 , n4282 , n310 );
    and g18916 ( n27061 , n11955 , n16894 );
    not g18917 ( n12189 , n31556 );
    and g18918 ( n8767 , n21101 , n27259 );
    nor g18919 ( n16034 , n29064 , n23723 );
    and g18920 ( n7117 , n23623 , n15067 );
    not g18921 ( n4895 , n13772 );
    not g18922 ( n27851 , n8085 );
    not g18923 ( n28500 , n20371 );
    xnor g18924 ( n15223 , n15221 , n18512 );
    nor g18925 ( n29151 , n18452 , n26306 );
    xnor g18926 ( n19776 , n3273 , n6705 );
    not g18927 ( n12335 , n29992 );
    not g18928 ( n14377 , n6534 );
    and g18929 ( n31374 , n3683 , n7297 );
    not g18930 ( n20546 , n1 );
    not g18931 ( n15666 , n25491 );
    xnor g18932 ( n14610 , n27042 , n7212 );
    xnor g18933 ( n25446 , n24350 , n24569 );
    xnor g18934 ( n1274 , n21136 , n9619 );
    xnor g18935 ( n14703 , n8453 , n16283 );
    nor g18936 ( n4208 , n20453 , n4623 );
    and g18937 ( n22275 , n6933 , n16351 );
    and g18938 ( n5253 , n8332 , n17296 );
    or g18939 ( n23945 , n19761 , n20223 );
    and g18940 ( n3183 , n30330 , n28813 );
    not g18941 ( n2820 , n11284 );
    not g18942 ( n939 , n17995 );
    and g18943 ( n30996 , n2724 , n9729 );
    xnor g18944 ( n3176 , n9840 , n19196 );
    not g18945 ( n4604 , n29253 );
    not g18946 ( n23459 , n20030 );
    not g18947 ( n24995 , n7270 );
    not g18948 ( n15582 , n4166 );
    not g18949 ( n10524 , n12264 );
    or g18950 ( n16965 , n10749 , n7078 );
    not g18951 ( n8961 , n7547 );
    nor g18952 ( n17706 , n7180 , n23651 );
    xnor g18953 ( n2382 , n31459 , n5170 );
    not g18954 ( n11050 , n9414 );
    and g18955 ( n16702 , n27439 , n9840 );
    not g18956 ( n8943 , n13924 );
    nor g18957 ( n4508 , n24525 , n10876 );
    or g18958 ( n249 , n25750 , n8973 );
    not g18959 ( n19444 , n7636 );
    xnor g18960 ( n16437 , n12803 , n14711 );
    and g18961 ( n7606 , n1034 , n31629 );
    xnor g18962 ( n10072 , n18439 , n17684 );
    not g18963 ( n16280 , n1275 );
    not g18964 ( n17493 , n14287 );
    and g18965 ( n12445 , n19829 , n23426 );
    xnor g18966 ( n16825 , n11973 , n14624 );
    and g18967 ( n17110 , n27164 , n27540 );
    or g18968 ( n2003 , n16675 , n20019 );
    not g18969 ( n23702 , n2186 );
    or g18970 ( n9493 , n17514 , n29584 );
    xnor g18971 ( n12032 , n3174 , n22941 );
    xnor g18972 ( n8161 , n17542 , n31294 );
    xnor g18973 ( n8267 , n15329 , n14641 );
    nor g18974 ( n15767 , n17499 , n9396 );
    not g18975 ( n15745 , n12160 );
    not g18976 ( n31638 , n17379 );
    not g18977 ( n3973 , n7323 );
    not g18978 ( n6123 , n13725 );
    or g18979 ( n16735 , n18389 , n13526 );
    or g18980 ( n10549 , n13948 , n21050 );
    and g18981 ( n19523 , n11455 , n25544 );
    xnor g18982 ( n3287 , n10476 , n7068 );
    or g18983 ( n24025 , n10484 , n7971 );
    nor g18984 ( n11465 , n14088 , n31750 );
    and g18985 ( n1101 , n27198 , n29492 );
    not g18986 ( n25597 , n24939 );
    not g18987 ( n21977 , n7471 );
    nor g18988 ( n20620 , n24614 , n30761 );
    nor g18989 ( n20336 , n7978 , n10316 );
    nor g18990 ( n11524 , n18025 , n19252 );
    or g18991 ( n13995 , n12148 , n31874 );
    or g18992 ( n15103 , n13468 , n10667 );
    and g18993 ( n10642 , n9051 , n20903 );
    or g18994 ( n4390 , n15567 , n24707 );
    and g18995 ( n21018 , n6241 , n12419 );
    and g18996 ( n31303 , n1821 , n1512 );
    and g18997 ( n26495 , n9275 , n4418 );
    or g18998 ( n9553 , n16953 , n10380 );
    and g18999 ( n21695 , n2208 , n8604 );
    not g19000 ( n11856 , n4973 );
    not g19001 ( n31401 , n19311 );
    not g19002 ( n22508 , n7591 );
    xnor g19003 ( n18224 , n30622 , n23703 );
    or g19004 ( n31269 , n2721 , n2967 );
    nor g19005 ( n2583 , n21464 , n23380 );
    not g19006 ( n4775 , n21049 );
    or g19007 ( n9576 , n24023 , n20923 );
    xnor g19008 ( n12908 , n29368 , n12803 );
    xnor g19009 ( n1337 , n1580 , n11331 );
    xnor g19010 ( n17005 , n7689 , n13763 );
    and g19011 ( n7758 , n29794 , n4924 );
    not g19012 ( n20940 , n8986 );
    and g19013 ( n1181 , n10858 , n1376 );
    and g19014 ( n441 , n4398 , n18157 );
    and g19015 ( n30599 , n24430 , n24629 );
    or g19016 ( n22201 , n8259 , n22714 );
    xnor g19017 ( n6993 , n29667 , n7651 );
    xor g19018 ( n10185 , n279 , n21809 );
    or g19019 ( n3112 , n7340 , n18564 );
    or g19020 ( n28476 , n24600 , n9724 );
    xnor g19021 ( n21577 , n10812 , n7241 );
    xnor g19022 ( n12988 , n26270 , n1717 );
    xnor g19023 ( n26698 , n16234 , n23764 );
    nor g19024 ( n4460 , n6217 , n2564 );
    or g19025 ( n7948 , n9139 , n17425 );
    xnor g19026 ( n17394 , n28081 , n14290 );
    xnor g19027 ( n20535 , n3155 , n18647 );
    not g19028 ( n30365 , n20431 );
    and g19029 ( n13844 , n8135 , n23225 );
    or g19030 ( n7372 , n2049 , n4934 );
    xnor g19031 ( n28024 , n30820 , n31489 );
    nor g19032 ( n21026 , n13495 , n2975 );
    or g19033 ( n12782 , n15507 , n2700 );
    nor g19034 ( n10213 , n138 , n29601 );
    xnor g19035 ( n10562 , n9248 , n481 );
    xnor g19036 ( n4990 , n490 , n7747 );
    xor g19037 ( n10978 , n31243 , n11461 );
    xnor g19038 ( n4073 , n8193 , n13457 );
    xnor g19039 ( n21970 , n5369 , n3423 );
    not g19040 ( n21130 , n10639 );
    not g19041 ( n8644 , n11838 );
    not g19042 ( n23882 , n16972 );
    xnor g19043 ( n18536 , n11609 , n13448 );
    not g19044 ( n16649 , n17262 );
    and g19045 ( n5430 , n24934 , n7697 );
    or g19046 ( n18261 , n7048 , n16430 );
    and g19047 ( n14111 , n15470 , n14180 );
    or g19048 ( n574 , n27719 , n14297 );
    and g19049 ( n11622 , n26575 , n13898 );
    and g19050 ( n15523 , n15965 , n2999 );
    not g19051 ( n11824 , n6704 );
    xnor g19052 ( n9005 , n11303 , n30887 );
    not g19053 ( n2357 , n23344 );
    or g19054 ( n18441 , n14729 , n18431 );
    and g19055 ( n22424 , n7058 , n20585 );
    or g19056 ( n4889 , n9000 , n7281 );
    nor g19057 ( n10074 , n7890 , n6738 );
    xnor g19058 ( n30336 , n24602 , n14066 );
    and g19059 ( n7941 , n28030 , n21843 );
    not g19060 ( n6118 , n4822 );
    and g19061 ( n4856 , n10294 , n15410 );
    not g19062 ( n26755 , n24607 );
    xnor g19063 ( n28822 , n11886 , n14356 );
    xnor g19064 ( n13846 , n27740 , n28951 );
    and g19065 ( n18482 , n432 , n25803 );
    or g19066 ( n11183 , n14144 , n20360 );
    or g19067 ( n12866 , n1254 , n5813 );
    and g19068 ( n765 , n1805 , n29916 );
    and g19069 ( n19214 , n2590 , n31612 );
    nor g19070 ( n16787 , n30046 , n16492 );
    xnor g19071 ( n17932 , n2400 , n20894 );
    or g19072 ( n28688 , n3447 , n20538 );
    xnor g19073 ( n10570 , n11984 , n28006 );
    not g19074 ( n29376 , n22521 );
    not g19075 ( n2976 , n5523 );
    xnor g19076 ( n3990 , n26754 , n16431 );
    or g19077 ( n14185 , n23419 , n21200 );
    not g19078 ( n13395 , n28884 );
    or g19079 ( n31967 , n13096 , n4303 );
    or g19080 ( n12005 , n10918 , n762 );
    xnor g19081 ( n14911 , n16970 , n6745 );
    or g19082 ( n9594 , n31355 , n5394 );
    or g19083 ( n15571 , n9496 , n8287 );
    and g19084 ( n8374 , n1092 , n21368 );
    not g19085 ( n12141 , n25414 );
    or g19086 ( n11496 , n1511 , n2266 );
    or g19087 ( n27377 , n5948 , n25958 );
    not g19088 ( n30992 , n6965 );
    not g19089 ( n13425 , n28170 );
    nor g19090 ( n1371 , n1084 , n23873 );
    or g19091 ( n26000 , n20946 , n12547 );
    and g19092 ( n23337 , n27231 , n27406 );
    nor g19093 ( n24831 , n25793 , n24137 );
    nor g19094 ( n11631 , n17617 , n10761 );
    and g19095 ( n30842 , n17922 , n28608 );
    or g19096 ( n12185 , n31974 , n21539 );
    xnor g19097 ( n24174 , n29367 , n1180 );
    or g19098 ( n25908 , n18548 , n2005 );
    not g19099 ( n10488 , n4326 );
    or g19100 ( n2696 , n14811 , n27105 );
    xnor g19101 ( n31266 , n11110 , n30562 );
    xnor g19102 ( n1064 , n6172 , n20510 );
    not g19103 ( n24280 , n30955 );
    not g19104 ( n1697 , n1997 );
    or g19105 ( n27879 , n7435 , n15024 );
    not g19106 ( n27511 , n28855 );
    not g19107 ( n12298 , n13701 );
    nor g19108 ( n23730 , n18667 , n8005 );
    or g19109 ( n20908 , n19910 , n14575 );
    xnor g19110 ( n405 , n26515 , n14745 );
    xnor g19111 ( n30906 , n6742 , n12566 );
    not g19112 ( n28211 , n9424 );
    not g19113 ( n21670 , n18274 );
    or g19114 ( n16458 , n20815 , n8994 );
    or g19115 ( n7067 , n3130 , n9899 );
    nor g19116 ( n31701 , n9595 , n16044 );
    or g19117 ( n1586 , n28871 , n16941 );
    and g19118 ( n12254 , n18231 , n31059 );
    nor g19119 ( n12348 , n16113 , n25904 );
    and g19120 ( n3107 , n8589 , n28459 );
    not g19121 ( n15080 , n24306 );
    and g19122 ( n9063 , n32 , n8468 );
    not g19123 ( n12527 , n2354 );
    and g19124 ( n13607 , n7086 , n23232 );
    xnor g19125 ( n5101 , n30450 , n18693 );
    xnor g19126 ( n23697 , n2005 , n26306 );
    or g19127 ( n22686 , n6034 , n31897 );
    xnor g19128 ( n2959 , n26445 , n15470 );
    not g19129 ( n1349 , n4451 );
    and g19130 ( n7302 , n1393 , n881 );
    xnor g19131 ( n5004 , n7283 , n6395 );
    or g19132 ( n13240 , n27791 , n29823 );
    nor g19133 ( n31129 , n10713 , n17584 );
    or g19134 ( n29969 , n17860 , n17900 );
    nor g19135 ( n16157 , n28350 , n26834 );
    not g19136 ( n10525 , n8764 );
    or g19137 ( n15553 , n31355 , n15668 );
    xnor g19138 ( n3326 , n14893 , n27413 );
    or g19139 ( n8591 , n20150 , n18662 );
    or g19140 ( n24293 , n31122 , n8805 );
    and g19141 ( n28378 , n13538 , n20965 );
    or g19142 ( n22112 , n3106 , n12098 );
    or g19143 ( n18745 , n20890 , n23801 );
    or g19144 ( n16460 , n30487 , n7289 );
    xnor g19145 ( n11306 , n27812 , n23310 );
    xnor g19146 ( n19466 , n3832 , n23779 );
    or g19147 ( n767 , n22887 , n10065 );
    or g19148 ( n26650 , n8523 , n24000 );
    not g19149 ( n331 , n24132 );
    not g19150 ( n24198 , n7254 );
    nor g19151 ( n28939 , n26349 , n31556 );
    or g19152 ( n9431 , n12777 , n27045 );
    or g19153 ( n25166 , n22039 , n2701 );
    not g19154 ( n7470 , n8839 );
    xnor g19155 ( n5079 , n5372 , n16178 );
    or g19156 ( n7441 , n21752 , n5162 );
    xnor g19157 ( n20397 , n23623 , n12256 );
    and g19158 ( n22529 , n26281 , n18378 );
    or g19159 ( n11780 , n7482 , n13857 );
    or g19160 ( n23302 , n23534 , n12292 );
    and g19161 ( n2901 , n22908 , n17804 );
    or g19162 ( n16770 , n27943 , n13942 );
    and g19163 ( n11751 , n20892 , n28295 );
    and g19164 ( n24261 , n4598 , n15910 );
    xnor g19165 ( n21502 , n13393 , n18165 );
    not g19166 ( n21441 , n28621 );
    or g19167 ( n30123 , n21176 , n3855 );
    and g19168 ( n16520 , n24270 , n14629 );
    not g19169 ( n13264 , n16861 );
    not g19170 ( n30104 , n14836 );
    xnor g19171 ( n22379 , n16818 , n6559 );
    nor g19172 ( n19532 , n788 , n4023 );
    not g19173 ( n2248 , n13526 );
    or g19174 ( n16907 , n23643 , n5215 );
    xnor g19175 ( n23299 , n16259 , n24712 );
    and g19176 ( n14302 , n12355 , n17090 );
    and g19177 ( n27790 , n20652 , n6195 );
    and g19178 ( n28539 , n28211 , n2825 );
    not g19179 ( n28238 , n24118 );
    nor g19180 ( n12750 , n25253 , n7644 );
    nor g19181 ( n16771 , n3755 , n13604 );
    xnor g19182 ( n18420 , n13942 , n30722 );
    nor g19183 ( n22410 , n20472 , n23138 );
    and g19184 ( n14080 , n16262 , n28966 );
    not g19185 ( n5532 , n22390 );
    not g19186 ( n41 , n23561 );
    xnor g19187 ( n11812 , n18824 , n10898 );
    not g19188 ( n27590 , n192 );
    xnor g19189 ( n17857 , n397 , n23934 );
    nor g19190 ( n11564 , n11850 , n8989 );
    not g19191 ( n22559 , n22941 );
    not g19192 ( n19929 , n19888 );
    xnor g19193 ( n27946 , n10246 , n18728 );
    xor g19194 ( n5194 , n21539 , n17371 );
    xnor g19195 ( n13644 , n29987 , n3948 );
    and g19196 ( n24077 , n23342 , n16803 );
    or g19197 ( n5009 , n28297 , n1687 );
    xnor g19198 ( n31205 , n9178 , n21531 );
    or g19199 ( n199 , n26670 , n9324 );
    not g19200 ( n28 , n11140 );
    not g19201 ( n14807 , n20326 );
    or g19202 ( n17545 , n2315 , n17771 );
    nor g19203 ( n762 , n3147 , n23593 );
    and g19204 ( n26744 , n19204 , n1732 );
    xnor g19205 ( n4384 , n31219 , n31998 );
    xnor g19206 ( n5670 , n6835 , n21873 );
    xor g19207 ( n24446 , n25779 , n23778 );
    xnor g19208 ( n7115 , n21943 , n19768 );
    xnor g19209 ( n16375 , n24290 , n5834 );
    xnor g19210 ( n14320 , n11554 , n15073 );
    or g19211 ( n2389 , n31499 , n9451 );
    or g19212 ( n9142 , n12030 , n6549 );
    xnor g19213 ( n29176 , n27432 , n31881 );
    not g19214 ( n1703 , n29186 );
    xnor g19215 ( n13914 , n30086 , n30969 );
    or g19216 ( n21065 , n21469 , n7588 );
    not g19217 ( n22934 , n16570 );
    not g19218 ( n4243 , n19801 );
    not g19219 ( n23369 , n13833 );
    xnor g19220 ( n14660 , n20807 , n6592 );
    or g19221 ( n21868 , n2200 , n6377 );
    xnor g19222 ( n1048 , n16849 , n2417 );
    not g19223 ( n23919 , n9270 );
    xnor g19224 ( n27985 , n10474 , n26114 );
    not g19225 ( n22806 , n31722 );
    not g19226 ( n9782 , n372 );
    xnor g19227 ( n1613 , n13402 , n8014 );
    not g19228 ( n19002 , n23094 );
    or g19229 ( n15605 , n21120 , n25383 );
    xnor g19230 ( n16201 , n24180 , n31910 );
    or g19231 ( n30626 , n10405 , n13159 );
    or g19232 ( n12545 , n6938 , n20839 );
    xnor g19233 ( n25778 , n5700 , n14583 );
    or g19234 ( n1558 , n18389 , n15424 );
    xnor g19235 ( n6872 , n8821 , n20351 );
    not g19236 ( n15022 , n2356 );
    not g19237 ( n28110 , n26203 );
    not g19238 ( n7344 , n21321 );
    not g19239 ( n31315 , n20057 );
    nor g19240 ( n21583 , n8529 , n28829 );
    and g19241 ( n12368 , n27691 , n29092 );
    and g19242 ( n18366 , n18897 , n12450 );
    nor g19243 ( n5044 , n15100 , n5864 );
    or g19244 ( n1904 , n15809 , n12822 );
    or g19245 ( n3263 , n5175 , n12720 );
    xor g19246 ( n26508 , n27232 , n30424 );
    not g19247 ( n1522 , n2329 );
    and g19248 ( n91 , n23434 , n2962 );
    not g19249 ( n15589 , n24522 );
    not g19250 ( n27006 , n26398 );
    not g19251 ( n31437 , n31539 );
    not g19252 ( n30387 , n15758 );
    or g19253 ( n6930 , n12558 , n15492 );
    not g19254 ( n8581 , n22776 );
    xnor g19255 ( n31202 , n10886 , n21104 );
    nor g19256 ( n29588 , n4532 , n22563 );
    nor g19257 ( n18146 , n28449 , n6111 );
    and g19258 ( n1940 , n18630 , n16781 );
    and g19259 ( n18757 , n16883 , n9161 );
    and g19260 ( n20268 , n25268 , n7178 );
    nor g19261 ( n18415 , n11132 , n23230 );
    or g19262 ( n12007 , n9920 , n2228 );
    not g19263 ( n27536 , n4484 );
    not g19264 ( n3057 , n24939 );
    and g19265 ( n14058 , n9513 , n16780 );
    nor g19266 ( n29264 , n2753 , n4258 );
    and g19267 ( n30410 , n14396 , n16066 );
    not g19268 ( n28366 , n7453 );
    or g19269 ( n29558 , n4166 , n510 );
    not g19270 ( n19802 , n13749 );
    not g19271 ( n4911 , n17162 );
    or g19272 ( n25225 , n20443 , n22693 );
    nor g19273 ( n20773 , n28058 , n3948 );
    and g19274 ( n13035 , n10194 , n3108 );
    nor g19275 ( n26407 , n18295 , n2932 );
    or g19276 ( n31793 , n29668 , n1841 );
    nor g19277 ( n25412 , n19570 , n20918 );
    nor g19278 ( n24962 , n624 , n28109 );
    xnor g19279 ( n24554 , n18789 , n5109 );
    xnor g19280 ( n22962 , n3112 , n28018 );
    not g19281 ( n3407 , n23839 );
    or g19282 ( n11335 , n1016 , n5571 );
    and g19283 ( n12240 , n28293 , n28517 );
    xnor g19284 ( n12804 , n30554 , n16461 );
    xnor g19285 ( n6407 , n21439 , n14786 );
    or g19286 ( n6718 , n2628 , n9235 );
    xnor g19287 ( n1434 , n9200 , n6046 );
    xnor g19288 ( n16937 , n18636 , n18352 );
    not g19289 ( n17638 , n21822 );
    or g19290 ( n12925 , n2108 , n21674 );
    not g19291 ( n13877 , n26676 );
    or g19292 ( n815 , n31292 , n18428 );
    not g19293 ( n11868 , n4376 );
    not g19294 ( n20519 , n22632 );
    and g19295 ( n6929 , n2881 , n28354 );
    xnor g19296 ( n9624 , n3641 , n7655 );
    or g19297 ( n9989 , n7457 , n1530 );
    xnor g19298 ( n25361 , n29764 , n25758 );
    xnor g19299 ( n21643 , n29731 , n12584 );
    or g19300 ( n30454 , n99 , n26925 );
    and g19301 ( n31174 , n21148 , n9640 );
    or g19302 ( n8746 , n13830 , n29464 );
    xnor g19303 ( n28767 , n17696 , n24835 );
    nor g19304 ( n3552 , n29519 , n9881 );
    or g19305 ( n26030 , n26551 , n2492 );
    not g19306 ( n26577 , n6295 );
    or g19307 ( n7339 , n28869 , n20267 );
    and g19308 ( n13403 , n15808 , n11967 );
    xnor g19309 ( n24187 , n8577 , n29252 );
    and g19310 ( n14455 , n20921 , n30900 );
    not g19311 ( n13614 , n21793 );
    xnor g19312 ( n29315 , n1266 , n9254 );
    xor g19313 ( n16655 , n14198 , n27591 );
    nor g19314 ( n13175 , n28381 , n20430 );
    not g19315 ( n24381 , n8134 );
    xnor g19316 ( n12220 , n19927 , n111 );
    and g19317 ( n23313 , n30373 , n17664 );
    or g19318 ( n7516 , n4142 , n9756 );
    xnor g19319 ( n5340 , n10099 , n31682 );
    not g19320 ( n23996 , n9693 );
    not g19321 ( n24517 , n7798 );
    xnor g19322 ( n26279 , n26039 , n10159 );
    or g19323 ( n22694 , n17414 , n27876 );
    not g19324 ( n19876 , n27926 );
    not g19325 ( n14999 , n18752 );
    or g19326 ( n6336 , n18596 , n29180 );
    nor g19327 ( n22510 , n20327 , n11655 );
    or g19328 ( n1001 , n11644 , n12773 );
    not g19329 ( n8803 , n2429 );
    xor g19330 ( n21362 , n15475 , n10149 );
    not g19331 ( n6377 , n12212 );
    and g19332 ( n680 , n14106 , n20262 );
    or g19333 ( n26403 , n18863 , n25576 );
    xnor g19334 ( n1218 , n9992 , n4833 );
    and g19335 ( n16753 , n25892 , n768 );
    or g19336 ( n8728 , n524 , n21449 );
    nor g19337 ( n31099 , n24512 , n30046 );
    and g19338 ( n29562 , n16754 , n19504 );
    xnor g19339 ( n13983 , n30731 , n9357 );
    and g19340 ( n23181 , n26184 , n16518 );
    not g19341 ( n26584 , n15878 );
    not g19342 ( n10909 , n30867 );
    nor g19343 ( n21853 , n7314 , n21374 );
    or g19344 ( n9296 , n2155 , n31410 );
    xnor g19345 ( n30393 , n4758 , n11619 );
    not g19346 ( n3997 , n6295 );
    not g19347 ( n28218 , n21767 );
    not g19348 ( n25902 , n3307 );
    not g19349 ( n9066 , n15672 );
    xnor g19350 ( n21089 , n13523 , n6810 );
    xnor g19351 ( n16869 , n23276 , n24225 );
    or g19352 ( n18618 , n5911 , n22636 );
    not g19353 ( n7545 , n4476 );
    and g19354 ( n13193 , n21905 , n7991 );
    or g19355 ( n24428 , n24831 , n3890 );
    not g19356 ( n22307 , n683 );
    xnor g19357 ( n23025 , n30314 , n20181 );
    not g19358 ( n24385 , n21595 );
    xnor g19359 ( n2202 , n8142 , n22453 );
    or g19360 ( n11160 , n22519 , n15323 );
    and g19361 ( n12523 , n9993 , n27103 );
    not g19362 ( n1863 , n30067 );
    xnor g19363 ( n11407 , n22288 , n27081 );
    xor g19364 ( n24391 , n2196 , n25353 );
    xnor g19365 ( n15774 , n7908 , n21311 );
    or g19366 ( n15420 , n3607 , n5179 );
    xnor g19367 ( n7532 , n3124 , n2818 );
    and g19368 ( n5278 , n28476 , n10575 );
    not g19369 ( n4815 , n11132 );
    or g19370 ( n25521 , n1986 , n11573 );
    xnor g19371 ( n3547 , n11943 , n30428 );
    or g19372 ( n27383 , n19577 , n23423 );
    not g19373 ( n32034 , n24493 );
    not g19374 ( n10907 , n4682 );
    xnor g19375 ( n1736 , n30382 , n8305 );
    not g19376 ( n22776 , n30427 );
    not g19377 ( n13840 , n7024 );
    or g19378 ( n27044 , n24018 , n2623 );
    not g19379 ( n19915 , n1449 );
    xnor g19380 ( n30124 , n24483 , n14271 );
    or g19381 ( n28753 , n13092 , n8782 );
    and g19382 ( n15713 , n29207 , n22664 );
    nor g19383 ( n22452 , n8550 , n27661 );
    and g19384 ( n31328 , n7197 , n12850 );
    or g19385 ( n9227 , n23991 , n17318 );
    not g19386 ( n28084 , n14477 );
    not g19387 ( n12673 , n22490 );
    or g19388 ( n31962 , n25037 , n8544 );
    not g19389 ( n12354 , n11381 );
    xor g19390 ( n27048 , n22241 , n23095 );
    nor g19391 ( n520 , n5948 , n13609 );
    xnor g19392 ( n17466 , n3821 , n1343 );
    and g19393 ( n30600 , n24563 , n4653 );
    xor g19394 ( n23779 , n31993 , n24939 );
    xnor g19395 ( n18010 , n20756 , n6527 );
    and g19396 ( n29526 , n29745 , n10676 );
    xnor g19397 ( n15544 , n14121 , n7009 );
    or g19398 ( n10178 , n30297 , n25851 );
    xnor g19399 ( n3157 , n29977 , n4089 );
    not g19400 ( n24824 , n5006 );
    and g19401 ( n21573 , n31541 , n10578 );
    nor g19402 ( n24715 , n30022 , n12815 );
    and g19403 ( n12276 , n24322 , n17796 );
    xnor g19404 ( n8235 , n3536 , n2921 );
    nor g19405 ( n6486 , n10543 , n22232 );
    xnor g19406 ( n31772 , n6955 , n8584 );
    or g19407 ( n12555 , n22803 , n13746 );
    nor g19408 ( n24816 , n24897 , n17236 );
    or g19409 ( n676 , n30794 , n13764 );
    not g19410 ( n11583 , n17001 );
    not g19411 ( n26783 , n9524 );
    not g19412 ( n7147 , n30529 );
    nor g19413 ( n20367 , n21122 , n21345 );
    or g19414 ( n29906 , n18394 , n13063 );
    xnor g19415 ( n29672 , n24191 , n14920 );
    not g19416 ( n8863 , n7937 );
    or g19417 ( n24168 , n18138 , n14152 );
    xnor g19418 ( n8380 , n29469 , n30113 );
    nor g19419 ( n12700 , n16524 , n7217 );
    and g19420 ( n12951 , n5659 , n30784 );
    and g19421 ( n30616 , n20858 , n27084 );
    nor g19422 ( n330 , n1985 , n4250 );
    and g19423 ( n424 , n22893 , n7953 );
    or g19424 ( n13223 , n17894 , n3572 );
    xnor g19425 ( n8090 , n26386 , n14516 );
    and g19426 ( n25070 , n10097 , n10389 );
    not g19427 ( n7128 , n29710 );
    or g19428 ( n21309 , n5331 , n16550 );
    or g19429 ( n2899 , n10435 , n25252 );
    xnor g19430 ( n17348 , n15834 , n687 );
    not g19431 ( n11271 , n8657 );
    not g19432 ( n6226 , n26266 );
    nor g19433 ( n23462 , n24725 , n8776 );
    xnor g19434 ( n29646 , n18328 , n15272 );
    not g19435 ( n26138 , n21358 );
    nor g19436 ( n15087 , n25838 , n26047 );
    or g19437 ( n26813 , n10959 , n24129 );
    xnor g19438 ( n13354 , n20999 , n1286 );
    or g19439 ( n17717 , n17839 , n22150 );
    nor g19440 ( n23217 , n13218 , n18254 );
    xnor g19441 ( n25398 , n14768 , n31639 );
    xnor g19442 ( n5778 , n10334 , n7046 );
    and g19443 ( n8556 , n27358 , n21213 );
    and g19444 ( n31640 , n8997 , n1969 );
    and g19445 ( n2888 , n17342 , n21272 );
    not g19446 ( n18443 , n23856 );
    xnor g19447 ( n13479 , n18038 , n19720 );
    not g19448 ( n26793 , n28462 );
    xnor g19449 ( n6358 , n4937 , n27185 );
    not g19450 ( n23890 , n14221 );
    or g19451 ( n19418 , n20601 , n11323 );
    xnor g19452 ( n9375 , n138 , n18391 );
    nor g19453 ( n10253 , n23556 , n2540 );
    nor g19454 ( n19745 , n8581 , n14843 );
    not g19455 ( n10373 , n16481 );
    and g19456 ( n153 , n2879 , n19848 );
    nor g19457 ( n15722 , n20519 , n21279 );
    or g19458 ( n31061 , n23110 , n9676 );
    buf g19459 ( n31414 , n12275 );
    nor g19460 ( n29944 , n24276 , n23666 );
    not g19461 ( n28766 , n11057 );
    not g19462 ( n2666 , n9812 );
    or g19463 ( n2867 , n4687 , n31400 );
    not g19464 ( n25599 , n13201 );
    and g19465 ( n24046 , n22153 , n15176 );
    nor g19466 ( n27877 , n18253 , n20599 );
    not g19467 ( n9714 , n25869 );
    not g19468 ( n4120 , n16301 );
    not g19469 ( n28282 , n3443 );
    nor g19470 ( n23220 , n5835 , n23458 );
    and g19471 ( n907 , n19486 , n2079 );
    xnor g19472 ( n21686 , n23569 , n28887 );
    or g19473 ( n23420 , n17833 , n29252 );
    not g19474 ( n15920 , n12335 );
    nor g19475 ( n11520 , n8245 , n24570 );
    not g19476 ( n15306 , n5683 );
    xor g19477 ( n19186 , n3247 , n9368 );
    xnor g19478 ( n12983 , n16232 , n29908 );
    nor g19479 ( n17161 , n1273 , n17437 );
    xnor g19480 ( n10054 , n20923 , n4335 );
    and g19481 ( n11691 , n21879 , n27455 );
    and g19482 ( n10651 , n13755 , n2481 );
    not g19483 ( n17279 , n9079 );
    or g19484 ( n7814 , n17406 , n29743 );
    and g19485 ( n20281 , n22365 , n17625 );
    and g19486 ( n3473 , n12157 , n29529 );
    xnor g19487 ( n8162 , n29818 , n4956 );
    nor g19488 ( n19382 , n23306 , n9653 );
    or g19489 ( n16898 , n14967 , n24304 );
    nor g19490 ( n11835 , n23115 , n1871 );
    not g19491 ( n2272 , n16856 );
    and g19492 ( n14568 , n22758 , n13044 );
    and g19493 ( n31510 , n31638 , n5243 );
    xnor g19494 ( n22643 , n19016 , n21076 );
    xnor g19495 ( n7671 , n163 , n21723 );
    nor g19496 ( n18047 , n12195 , n5545 );
    not g19497 ( n22598 , n1633 );
    xnor g19498 ( n21796 , n26200 , n29180 );
    xnor g19499 ( n26218 , n18517 , n29252 );
    nor g19500 ( n29723 , n10034 , n30505 );
    and g19501 ( n30963 , n18805 , n13042 );
    nor g19502 ( n17564 , n17887 , n22361 );
    and g19503 ( n22780 , n1843 , n16020 );
    not g19504 ( n5864 , n23744 );
    or g19505 ( n18535 , n9411 , n11764 );
    buf g19506 ( n4701 , n29932 );
    and g19507 ( n21195 , n6827 , n10792 );
    xnor g19508 ( n26251 , n29764 , n21122 );
    or g19509 ( n23831 , n14096 , n3972 );
    nor g19510 ( n976 , n28776 , n25986 );
    xnor g19511 ( n29697 , n28417 , n6888 );
    or g19512 ( n29775 , n14686 , n10607 );
    not g19513 ( n23287 , n24758 );
    nor g19514 ( n25079 , n20597 , n16461 );
    or g19515 ( n25983 , n15147 , n22428 );
    and g19516 ( n29876 , n8748 , n31146 );
    and g19517 ( n11417 , n14933 , n18173 );
    not g19518 ( n11166 , n3076 );
    not g19519 ( n4723 , n30067 );
    xnor g19520 ( n13562 , n27446 , n7990 );
    not g19521 ( n9859 , n10759 );
    and g19522 ( n1338 , n14429 , n1245 );
    not g19523 ( n18537 , n17651 );
    nor g19524 ( n26951 , n6859 , n26561 );
    xnor g19525 ( n21298 , n9948 , n16238 );
    and g19526 ( n28017 , n13297 , n4035 );
    not g19527 ( n21326 , n11716 );
    nor g19528 ( n21043 , n6527 , n11601 );
    or g19529 ( n13143 , n13410 , n11649 );
    or g19530 ( n30066 , n29437 , n679 );
    nor g19531 ( n2827 , n5456 , n15778 );
    not g19532 ( n12182 , n4145 );
    xnor g19533 ( n15449 , n3175 , n15745 );
    xnor g19534 ( n18608 , n2519 , n31603 );
    xnor g19535 ( n7188 , n16815 , n6603 );
    nor g19536 ( n28416 , n24216 , n23217 );
    not g19537 ( n12774 , n5544 );
    xnor g19538 ( n19911 , n18647 , n7787 );
    or g19539 ( n15114 , n1407 , n1243 );
    and g19540 ( n23333 , n15926 , n12008 );
    or g19541 ( n19154 , n21847 , n22083 );
    xnor g19542 ( n21223 , n19255 , n4836 );
    xnor g19543 ( n31372 , n19948 , n9205 );
    and g19544 ( n19626 , n4387 , n11437 );
    nor g19545 ( n11201 , n1915 , n1471 );
    xnor g19546 ( n17947 , n27775 , n27359 );
    not g19547 ( n11439 , n30616 );
    not g19548 ( n24402 , n23071 );
    xnor g19549 ( n24564 , n2296 , n27896 );
    or g19550 ( n10536 , n11584 , n31809 );
    and g19551 ( n15490 , n9041 , n10877 );
    xnor g19552 ( n17505 , n20156 , n23023 );
    and g19553 ( n26288 , n9207 , n10896 );
    xnor g19554 ( n30830 , n10307 , n23013 );
    xnor g19555 ( n9590 , n19069 , n22606 );
    not g19556 ( n19248 , n29239 );
    xnor g19557 ( n27832 , n23907 , n29444 );
    xnor g19558 ( n22232 , n21586 , n8428 );
    and g19559 ( n1963 , n15242 , n21281 );
    and g19560 ( n11080 , n10150 , n11466 );
    or g19561 ( n5177 , n31120 , n31375 );
    or g19562 ( n24650 , n29401 , n27817 );
    xnor g19563 ( n15464 , n29764 , n4662 );
    xnor g19564 ( n22350 , n23257 , n8561 );
    or g19565 ( n15244 , n9389 , n6085 );
    and g19566 ( n10091 , n24732 , n3655 );
    xnor g19567 ( n4953 , n4859 , n17851 );
    nor g19568 ( n8905 , n2683 , n4730 );
    not g19569 ( n17796 , n24913 );
    not g19570 ( n2139 , n23277 );
    not g19571 ( n17325 , n30340 );
    or g19572 ( n27989 , n1351 , n11669 );
    or g19573 ( n17964 , n4947 , n29946 );
    xnor g19574 ( n30845 , n16 , n23962 );
    xnor g19575 ( n10626 , n20471 , n18612 );
    xnor g19576 ( n8854 , n12519 , n13939 );
    xnor g19577 ( n17855 , n4251 , n6934 );
    xnor g19578 ( n824 , n27198 , n4555 );
    not g19579 ( n1861 , n13262 );
    not g19580 ( n3118 , n23137 );
    or g19581 ( n27076 , n3440 , n10669 );
    not g19582 ( n73 , n14555 );
    not g19583 ( n22576 , n13813 );
    not g19584 ( n10787 , n4844 );
    or g19585 ( n23586 , n30002 , n26894 );
    nor g19586 ( n529 , n16209 , n28638 );
    and g19587 ( n8938 , n26459 , n17138 );
    not g19588 ( n29079 , n13955 );
    xnor g19589 ( n5345 , n3561 , n18432 );
    not g19590 ( n12277 , n16462 );
    nor g19591 ( n8329 , n9136 , n21986 );
    not g19592 ( n6721 , n15292 );
    not g19593 ( n8056 , n26934 );
    or g19594 ( n15757 , n24319 , n29979 );
    not g19595 ( n2606 , n5166 );
    xnor g19596 ( n24416 , n13569 , n19153 );
    xnor g19597 ( n31294 , n13442 , n1738 );
    not g19598 ( n20456 , n1461 );
    xnor g19599 ( n4472 , n8233 , n23886 );
    or g19600 ( n26141 , n12124 , n22779 );
    and g19601 ( n16698 , n15832 , n25540 );
    not g19602 ( n353 , n23226 );
    and g19603 ( n21539 , n26263 , n25224 );
    not g19604 ( n17959 , n3251 );
    not g19605 ( n10332 , n6216 );
    or g19606 ( n5516 , n20548 , n20602 );
    xnor g19607 ( n8221 , n8814 , n4132 );
    not g19608 ( n10861 , n27487 );
    or g19609 ( n16949 , n22549 , n731 );
    not g19610 ( n23833 , n29834 );
    xnor g19611 ( n27449 , n27829 , n14503 );
    not g19612 ( n26473 , n15195 );
    or g19613 ( n31418 , n5629 , n8817 );
    xnor g19614 ( n10561 , n25669 , n25006 );
    not g19615 ( n30519 , n20825 );
    xnor g19616 ( n25813 , n29540 , n13800 );
    or g19617 ( n17942 , n9382 , n10585 );
    or g19618 ( n8395 , n937 , n2734 );
    xnor g19619 ( n24325 , n23161 , n10250 );
    or g19620 ( n4537 , n18325 , n18581 );
    or g19621 ( n10702 , n16446 , n22459 );
    xnor g19622 ( n26186 , n5970 , n5662 );
    not g19623 ( n11608 , n9011 );
    or g19624 ( n15697 , n289 , n7929 );
    not g19625 ( n24697 , n31246 );
    xnor g19626 ( n4530 , n14606 , n24456 );
    or g19627 ( n11483 , n21534 , n2378 );
    xnor g19628 ( n4698 , n28096 , n5077 );
    xnor g19629 ( n10075 , n29479 , n17929 );
    not g19630 ( n9973 , n19080 );
    or g19631 ( n27932 , n30471 , n25176 );
    not g19632 ( n6246 , n11643 );
    or g19633 ( n32023 , n7822 , n25615 );
    not g19634 ( n29338 , n188 );
    and g19635 ( n13455 , n5669 , n21978 );
    or g19636 ( n631 , n26636 , n12779 );
    and g19637 ( n17182 , n1878 , n13383 );
    nor g19638 ( n27560 , n5388 , n17854 );
    nor g19639 ( n32014 , n2001 , n6058 );
    or g19640 ( n10465 , n19809 , n17988 );
    and g19641 ( n1449 , n24997 , n8011 );
    or g19642 ( n841 , n25279 , n5163 );
    and g19643 ( n6772 , n5714 , n11558 );
    or g19644 ( n14355 , n18696 , n4107 );
    xnor g19645 ( n5733 , n6714 , n6306 );
    or g19646 ( n23672 , n2706 , n5630 );
    nor g19647 ( n19757 , n25599 , n22637 );
    not g19648 ( n1025 , n4159 );
    not g19649 ( n16804 , n11469 );
    not g19650 ( n3544 , n25730 );
    nor g19651 ( n18883 , n31895 , n10005 );
    and g19652 ( n26831 , n8712 , n24807 );
    or g19653 ( n27984 , n20632 , n13393 );
    xnor g19654 ( n21409 , n1957 , n28180 );
    not g19655 ( n10936 , n15582 );
    or g19656 ( n27281 , n4812 , n20318 );
    not g19657 ( n6429 , n11218 );
    not g19658 ( n31250 , n20526 );
    or g19659 ( n10694 , n11298 , n27031 );
    or g19660 ( n7189 , n15216 , n20377 );
    xnor g19661 ( n23174 , n19802 , n24387 );
    nor g19662 ( n496 , n19425 , n1997 );
    or g19663 ( n23079 , n15533 , n31149 );
    xor g19664 ( n13672 , n9404 , n1127 );
    xnor g19665 ( n29417 , n27376 , n17159 );
    not g19666 ( n27207 , n31989 );
    and g19667 ( n31509 , n18079 , n18663 );
    and g19668 ( n26515 , n17383 , n11186 );
    not g19669 ( n21258 , n17617 );
    xnor g19670 ( n8733 , n4036 , n13135 );
    or g19671 ( n30109 , n15261 , n24247 );
    and g19672 ( n30890 , n23067 , n3210 );
    xnor g19673 ( n246 , n13868 , n10574 );
    xnor g19674 ( n740 , n10720 , n1628 );
    or g19675 ( n16988 , n7013 , n26585 );
    or g19676 ( n27110 , n23044 , n353 );
    xnor g19677 ( n1773 , n25913 , n16019 );
    and g19678 ( n22533 , n31178 , n16728 );
    or g19679 ( n20353 , n8000 , n3720 );
    nor g19680 ( n20395 , n10521 , n4608 );
    or g19681 ( n4806 , n11736 , n675 );
    buf g19682 ( n20630 , n25462 );
    nor g19683 ( n4110 , n6639 , n29664 );
    or g19684 ( n9422 , n27398 , n22987 );
    xnor g19685 ( n26467 , n29422 , n27964 );
    and g19686 ( n15153 , n17435 , n16598 );
    not g19687 ( n25668 , n18253 );
    and g19688 ( n4272 , n15272 , n1736 );
    not g19689 ( n28394 , n3907 );
    xnor g19690 ( n22096 , n7277 , n28433 );
    or g19691 ( n17061 , n26114 , n26066 );
    xnor g19692 ( n22946 , n30447 , n13209 );
    not g19693 ( n24023 , n28433 );
    nor g19694 ( n10867 , n1720 , n21185 );
    or g19695 ( n27102 , n25338 , n13549 );
    nor g19696 ( n9451 , n10806 , n16167 );
    xnor g19697 ( n827 , n2383 , n19256 );
    xnor g19698 ( n3773 , n30935 , n8872 );
    or g19699 ( n27823 , n7960 , n2415 );
    or g19700 ( n5785 , n11291 , n11968 );
    or g19701 ( n860 , n5368 , n7695 );
    xnor g19702 ( n9772 , n12478 , n18394 );
    not g19703 ( n21153 , n21454 );
    or g19704 ( n17088 , n6177 , n20910 );
    not g19705 ( n7753 , n19710 );
    not g19706 ( n8289 , n19262 );
    nor g19707 ( n849 , n20994 , n15245 );
    not g19708 ( n23026 , n11440 );
    xnor g19709 ( n21949 , n19425 , n1997 );
    not g19710 ( n16333 , n28319 );
    nor g19711 ( n27656 , n4451 , n11157 );
    and g19712 ( n15549 , n2000 , n17019 );
    not g19713 ( n8023 , n30923 );
    not g19714 ( n299 , n7742 );
    nor g19715 ( n8209 , n24985 , n11603 );
    or g19716 ( n11842 , n15138 , n16527 );
    not g19717 ( n11391 , n30557 );
    not g19718 ( n14950 , n18474 );
    or g19719 ( n5335 , n14457 , n3998 );
    not g19720 ( n4978 , n17753 );
    or g19721 ( n7783 , n26529 , n6280 );
    xnor g19722 ( n4160 , n10756 , n30643 );
    or g19723 ( n11358 , n27878 , n3143 );
    or g19724 ( n23152 , n2103 , n31671 );
    not g19725 ( n18114 , n19241 );
    not g19726 ( n16763 , n15792 );
    xor g19727 ( n6591 , n10487 , n4804 );
    or g19728 ( n23384 , n8608 , n14482 );
    xnor g19729 ( n31134 , n23782 , n3411 );
    not g19730 ( n8474 , n10477 );
    xnor g19731 ( n12733 , n7542 , n17617 );
    or g19732 ( n26238 , n287 , n9857 );
    and g19733 ( n86 , n25851 , n30297 );
    xnor g19734 ( n6388 , n17344 , n7235 );
    not g19735 ( n8364 , n2457 );
    xnor g19736 ( n589 , n25301 , n3990 );
    not g19737 ( n21902 , n2971 );
    or g19738 ( n5303 , n1035 , n3975 );
    not g19739 ( n1288 , n7839 );
    nor g19740 ( n3542 , n24988 , n27906 );
    xnor g19741 ( n19229 , n11622 , n16359 );
    nor g19742 ( n14549 , n12306 , n20005 );
    xor g19743 ( n16410 , n29625 , n29041 );
    not g19744 ( n11721 , n28252 );
    xnor g19745 ( n27741 , n29328 , n29725 );
    not g19746 ( n8163 , n9043 );
    xnor g19747 ( n18865 , n515 , n13549 );
    xnor g19748 ( n27602 , n6241 , n14988 );
    not g19749 ( n15158 , n17325 );
    and g19750 ( n24846 , n284 , n635 );
    and g19751 ( n5865 , n5878 , n30538 );
    nor g19752 ( n25161 , n8714 , n2248 );
    nor g19753 ( n27489 , n20041 , n23995 );
    or g19754 ( n20004 , n443 , n21079 );
    xnor g19755 ( n3488 , n4088 , n7310 );
    not g19756 ( n23926 , n28616 );
    or g19757 ( n14725 , n19215 , n5028 );
    not g19758 ( n16109 , n614 );
    buf g19759 ( n31355 , n30957 );
    xnor g19760 ( n19056 , n1248 , n3094 );
    xnor g19761 ( n30141 , n8646 , n7926 );
    not g19762 ( n12754 , n29471 );
    not g19763 ( n25218 , n21350 );
    buf g19764 ( n19282 , n31566 );
    and g19765 ( n1949 , n16305 , n11376 );
    and g19766 ( n5128 , n28789 , n13980 );
    xnor g19767 ( n2420 , n1675 , n9336 );
    not g19768 ( n18852 , n10028 );
    or g19769 ( n12906 , n25650 , n6772 );
    xnor g19770 ( n14345 , n11172 , n29321 );
    xnor g19771 ( n5949 , n23260 , n3579 );
    not g19772 ( n27169 , n27946 );
    and g19773 ( n17345 , n17433 , n8916 );
    nor g19774 ( n20062 , n28238 , n6917 );
    and g19775 ( n13058 , n28346 , n2060 );
    and g19776 ( n20079 , n29150 , n26165 );
    or g19777 ( n2480 , n28968 , n6280 );
    not g19778 ( n10252 , n22574 );
    nor g19779 ( n23642 , n27309 , n20456 );
    not g19780 ( n20408 , n27086 );
    xnor g19781 ( n22690 , n20809 , n24652 );
    not g19782 ( n13647 , n12384 );
    xor g19783 ( n12201 , n12139 , n19466 );
    xnor g19784 ( n1679 , n26605 , n8082 );
    xnor g19785 ( n7007 , n25808 , n5131 );
    not g19786 ( n20597 , n28588 );
    not g19787 ( n5312 , n29643 );
    not g19788 ( n1044 , n30396 );
    and g19789 ( n9965 , n18635 , n25775 );
    not g19790 ( n12688 , n2723 );
    not g19791 ( n20123 , n9901 );
    not g19792 ( n13553 , n23919 );
    or g19793 ( n8656 , n2937 , n25798 );
    xor g19794 ( n2937 , n10085 , n14379 );
    nor g19795 ( n31611 , n19340 , n5133 );
    xnor g19796 ( n1699 , n8465 , n2069 );
    xnor g19797 ( n535 , n28065 , n13698 );
    or g19798 ( n26124 , n29768 , n20734 );
    nor g19799 ( n28007 , n17764 , n17614 );
    xnor g19800 ( n1405 , n23195 , n10433 );
    not g19801 ( n494 , n1281 );
    xnor g19802 ( n3605 , n31896 , n30525 );
    and g19803 ( n12848 , n6821 , n27191 );
    and g19804 ( n23909 , n6731 , n9682 );
    nor g19805 ( n31056 , n19055 , n12498 );
    not g19806 ( n27957 , n15055 );
    or g19807 ( n24329 , n7124 , n886 );
    nor g19808 ( n30924 , n15993 , n19183 );
    xnor g19809 ( n24940 , n14407 , n3775 );
    and g19810 ( n7726 , n3913 , n6170 );
    xnor g19811 ( n6818 , n25377 , n31614 );
    and g19812 ( n24798 , n4308 , n6119 );
    or g19813 ( n25885 , n4576 , n2823 );
    xnor g19814 ( n31189 , n39 , n13521 );
    not g19815 ( n20913 , n5071 );
    not g19816 ( n2283 , n21911 );
    not g19817 ( n30917 , n11905 );
    not g19818 ( n17204 , n3614 );
    not g19819 ( n25179 , n25037 );
    not g19820 ( n29142 , n3361 );
    not g19821 ( n5923 , n16719 );
    xnor g19822 ( n808 , n21401 , n7898 );
    or g19823 ( n31321 , n22212 , n10244 );
    nor g19824 ( n20568 , n27682 , n2220 );
    nor g19825 ( n18602 , n20905 , n21925 );
    xnor g19826 ( n9067 , n27614 , n28404 );
    not g19827 ( n21047 , n9830 );
    xnor g19828 ( n29462 , n1303 , n12911 );
    and g19829 ( n18703 , n18740 , n10039 );
    not g19830 ( n25182 , n18065 );
    not g19831 ( n28202 , n4451 );
    and g19832 ( n29690 , n7449 , n17361 );
    or g19833 ( n28595 , n25515 , n351 );
    not g19834 ( n8225 , n29075 );
    and g19835 ( n602 , n31663 , n11556 );
    and g19836 ( n2585 , n25942 , n31468 );
    and g19837 ( n21759 , n2719 , n20664 );
    or g19838 ( n28553 , n21060 , n17700 );
    and g19839 ( n11503 , n23073 , n26057 );
    or g19840 ( n16009 , n9043 , n9163 );
    or g19841 ( n5859 , n26420 , n6339 );
    and g19842 ( n12300 , n24332 , n1776 );
    and g19843 ( n31358 , n3833 , n10535 );
    or g19844 ( n28485 , n4906 , n13506 );
    xnor g19845 ( n20338 , n28244 , n28019 );
    not g19846 ( n23954 , n28734 );
    xnor g19847 ( n27958 , n4581 , n6977 );
    or g19848 ( n29572 , n11142 , n27629 );
    not g19849 ( n5845 , n7144 );
    xor g19850 ( n6925 , n855 , n31102 );
    not g19851 ( n6352 , n8806 );
    or g19852 ( n31530 , n9928 , n11510 );
    xnor g19853 ( n6612 , n30392 , n16879 );
    xnor g19854 ( n7641 , n23668 , n7190 );
    or g19855 ( n20061 , n11051 , n8874 );
    or g19856 ( n31630 , n15761 , n17369 );
    or g19857 ( n3827 , n5260 , n19892 );
    not g19858 ( n7152 , n19721 );
    or g19859 ( n11158 , n24739 , n20695 );
    not g19860 ( n15439 , n17895 );
    and g19861 ( n27251 , n31039 , n4062 );
    or g19862 ( n30116 , n21926 , n4339 );
    and g19863 ( n6786 , n15493 , n20304 );
    not g19864 ( n30062 , n28009 );
    not g19865 ( n18470 , n26591 );
    and g19866 ( n8528 , n11765 , n12024 );
    xnor g19867 ( n2397 , n2924 , n2665 );
    or g19868 ( n23874 , n23896 , n25390 );
    or g19869 ( n25054 , n11254 , n18014 );
    xor g19870 ( n17790 , n26347 , n420 );
    or g19871 ( n30081 , n13568 , n24266 );
    not g19872 ( n4802 , n27589 );
    and g19873 ( n26832 , n19252 , n18025 );
    and g19874 ( n24426 , n11030 , n10219 );
    not g19875 ( n11175 , n28288 );
    and g19876 ( n6884 , n13361 , n889 );
    not g19877 ( n28226 , n4480 );
    not g19878 ( n12684 , n11618 );
    and g19879 ( n2155 , n14290 , n23852 );
    or g19880 ( n8448 , n2386 , n948 );
    and g19881 ( n26180 , n623 , n20520 );
    xnor g19882 ( n1880 , n17434 , n6577 );
    not g19883 ( n12863 , n22670 );
    xnor g19884 ( n10728 , n14334 , n19421 );
    xnor g19885 ( n17054 , n20279 , n15830 );
    nor g19886 ( n18225 , n3108 , n14377 );
    not g19887 ( n31231 , n20339 );
    or g19888 ( n10849 , n20833 , n28101 );
    or g19889 ( n10392 , n10144 , n11686 );
    not g19890 ( n18840 , n654 );
    not g19891 ( n15221 , n12211 );
    or g19892 ( n27358 , n12168 , n25528 );
    not g19893 ( n12309 , n11792 );
    and g19894 ( n8708 , n522 , n11843 );
    not g19895 ( n4827 , n28845 );
    not g19896 ( n10946 , n22573 );
    xnor g19897 ( n21300 , n8030 , n21960 );
    and g19898 ( n28171 , n14263 , n7581 );
    not g19899 ( n28134 , n21760 );
    xnor g19900 ( n16228 , n12179 , n6507 );
    xnor g19901 ( n25945 , n22070 , n10974 );
    not g19902 ( n10210 , n1678 );
    xor g19903 ( n10129 , n19953 , n24344 );
    nor g19904 ( n19419 , n204 , n23652 );
    xnor g19905 ( n29054 , n15382 , n26598 );
    xnor g19906 ( n3323 , n14459 , n8143 );
    and g19907 ( n7530 , n24051 , n24904 );
    xnor g19908 ( n24194 , n19211 , n27355 );
    xnor g19909 ( n20837 , n10878 , n31937 );
    xnor g19910 ( n13363 , n3673 , n10113 );
    and g19911 ( n31717 , n17717 , n19018 );
    xnor g19912 ( n23757 , n4233 , n13621 );
    not g19913 ( n4347 , n2331 );
    xnor g19914 ( n4132 , n1616 , n30405 );
    nor g19915 ( n14865 , n8423 , n150 );
    xnor g19916 ( n18519 , n14562 , n14707 );
    or g19917 ( n27445 , n13087 , n15524 );
    not g19918 ( n12443 , n8988 );
    and g19919 ( n28041 , n7877 , n24094 );
    or g19920 ( n2094 , n9744 , n19892 );
    not g19921 ( n20101 , n19295 );
    not g19922 ( n15730 , n25360 );
    and g19923 ( n13214 , n6762 , n19828 );
    not g19924 ( n9924 , n22395 );
    not g19925 ( n20435 , n15772 );
    xnor g19926 ( n16518 , n2896 , n1892 );
    and g19927 ( n22993 , n26215 , n13163 );
    or g19928 ( n31663 , n5787 , n14647 );
    and g19929 ( n19040 , n22229 , n19515 );
    and g19930 ( n20477 , n12886 , n21423 );
    and g19931 ( n19113 , n28919 , n17227 );
    not g19932 ( n21135 , n9582 );
    not g19933 ( n28207 , n26969 );
    or g19934 ( n28970 , n19489 , n15470 );
    and g19935 ( n31256 , n5920 , n18314 );
    not g19936 ( n6701 , n20894 );
    not g19937 ( n12849 , n16115 );
    xnor g19938 ( n3285 , n7929 , n16271 );
    and g19939 ( n29043 , n3231 , n18952 );
    xor g19940 ( n17900 , n441 , n21603 );
    or g19941 ( n25604 , n27701 , n4802 );
    xnor g19942 ( n16166 , n25324 , n7068 );
    or g19943 ( n12465 , n20390 , n11667 );
    xnor g19944 ( n22713 , n3227 , n7730 );
    not g19945 ( n20680 , n8964 );
    not g19946 ( n12013 , n14361 );
    xnor g19947 ( n5725 , n21104 , n4257 );
    nor g19948 ( n4919 , n28672 , n16353 );
    xnor g19949 ( n28713 , n4701 , n17149 );
    not g19950 ( n18837 , n15074 );
    and g19951 ( n30627 , n14964 , n8581 );
    or g19952 ( n14120 , n25692 , n18172 );
    xnor g19953 ( n26075 , n20412 , n27501 );
    nor g19954 ( n31952 , n28546 , n29796 );
    and g19955 ( n5990 , n22380 , n31279 );
    xnor g19956 ( n27754 , n21136 , n19217 );
    xnor g19957 ( n23572 , n5918 , n10846 );
    or g19958 ( n27188 , n3615 , n30582 );
    not g19959 ( n17597 , n10696 );
    not g19960 ( n2855 , n16604 );
    xnor g19961 ( n7345 , n13481 , n7455 );
    and g19962 ( n3071 , n23466 , n870 );
    buf g19963 ( n2704 , n24901 );
    not g19964 ( n11484 , n9374 );
    and g19965 ( n25102 , n9388 , n18082 );
    xnor g19966 ( n6200 , n4598 , n11349 );
    and g19967 ( n3674 , n12643 , n14404 );
    xnor g19968 ( n9582 , n4094 , n20242 );
    or g19969 ( n16065 , n2153 , n4212 );
    and g19970 ( n17169 , n14643 , n15009 );
    or g19971 ( n16902 , n1977 , n10841 );
    xnor g19972 ( n6632 , n10351 , n19596 );
    not g19973 ( n11392 , n5262 );
    nor g19974 ( n23243 , n24366 , n15950 );
    and g19975 ( n21828 , n10087 , n27945 );
    or g19976 ( n14497 , n20135 , n27820 );
    and g19977 ( n18790 , n12382 , n29969 );
    not g19978 ( n4037 , n23510 );
    xnor g19979 ( n5192 , n2246 , n20872 );
    and g19980 ( n9407 , n1082 , n5896 );
    xnor g19981 ( n30105 , n3126 , n20662 );
    xnor g19982 ( n1579 , n8701 , n8921 );
    and g19983 ( n18614 , n14275 , n4506 );
    not g19984 ( n24308 , n14536 );
    xnor g19985 ( n29234 , n4216 , n22350 );
    not g19986 ( n12929 , n8520 );
    or g19987 ( n19321 , n7068 , n449 );
    not g19988 ( n3869 , n16845 );
    nor g19989 ( n22892 , n5625 , n9156 );
    xnor g19990 ( n29375 , n8866 , n21866 );
    and g19991 ( n31601 , n4433 , n23017 );
    or g19992 ( n26617 , n8063 , n4072 );
    xnor g19993 ( n12481 , n25276 , n26758 );
    or g19994 ( n22000 , n242 , n29469 );
    xnor g19995 ( n4013 , n7209 , n27453 );
    not g19996 ( n27115 , n12212 );
    xnor g19997 ( n5806 , n26332 , n7014 );
    and g19998 ( n16857 , n20972 , n2361 );
    xnor g19999 ( n30577 , n29069 , n29439 );
    or g20000 ( n27595 , n30457 , n9589 );
    or g20001 ( n9421 , n1650 , n18848 );
    and g20002 ( n21346 , n1354 , n9495 );
    xor g20003 ( n19057 , n2383 , n17954 );
    and g20004 ( n3497 , n25050 , n24065 );
    not g20005 ( n6404 , n6872 );
    and g20006 ( n31691 , n11481 , n12318 );
    not g20007 ( n7452 , n15636 );
    nor g20008 ( n3349 , n27002 , n30607 );
    not g20009 ( n6661 , n23172 );
    nor g20010 ( n6248 , n9345 , n8285 );
    xnor g20011 ( n24452 , n12851 , n10606 );
    xnor g20012 ( n6477 , n28892 , n13393 );
    xnor g20013 ( n12827 , n3371 , n8419 );
    or g20014 ( n14873 , n26306 , n20680 );
    or g20015 ( n15371 , n20612 , n2285 );
    not g20016 ( n13576 , n25397 );
    xnor g20017 ( n18995 , n426 , n17646 );
    and g20018 ( n30223 , n1174 , n28595 );
    not g20019 ( n20438 , n11574 );
    nor g20020 ( n30612 , n3345 , n22631 );
    and g20021 ( n14429 , n10686 , n28239 );
    xnor g20022 ( n15226 , n28707 , n20052 );
    or g20023 ( n21576 , n4348 , n22859 );
    xnor g20024 ( n30999 , n21092 , n1637 );
    or g20025 ( n19318 , n24024 , n24982 );
    not g20026 ( n20850 , n17317 );
    xnor g20027 ( n3433 , n23065 , n17348 );
    not g20028 ( n19845 , n30706 );
    and g20029 ( n16539 , n24623 , n26416 );
    not g20030 ( n4086 , n27101 );
    not g20031 ( n20515 , n831 );
    or g20032 ( n18365 , n16356 , n6152 );
    not g20033 ( n24396 , n19590 );
    xnor g20034 ( n20636 , n14555 , n9591 );
    nor g20035 ( n16032 , n590 , n3616 );
    not g20036 ( n7377 , n21261 );
    xnor g20037 ( n4764 , n9923 , n9113 );
    not g20038 ( n17595 , n21846 );
    and g20039 ( n1061 , n1753 , n8113 );
    not g20040 ( n10828 , n2054 );
    nor g20041 ( n1386 , n8352 , n411 );
    nor g20042 ( n12932 , n4875 , n30865 );
    and g20043 ( n19487 , n15378 , n31162 );
    not g20044 ( n28012 , n29702 );
    xnor g20045 ( n16841 , n9424 , n9653 );
    xnor g20046 ( n30213 , n31783 , n21508 );
    xnor g20047 ( n23335 , n20757 , n11956 );
    not g20048 ( n29780 , n10411 );
    and g20049 ( n26806 , n7618 , n27460 );
    or g20050 ( n6918 , n11172 , n30898 );
    and g20051 ( n24958 , n21 , n31891 );
    and g20052 ( n16085 , n2068 , n31908 );
    and g20053 ( n17370 , n22311 , n28668 );
    xnor g20054 ( n19333 , n18625 , n776 );
    not g20055 ( n12940 , n6040 );
    and g20056 ( n4683 , n9715 , n11652 );
    xnor g20057 ( n10350 , n8135 , n14383 );
    not g20058 ( n14499 , n22045 );
    or g20059 ( n26402 , n4061 , n24898 );
    and g20060 ( n28923 , n22186 , n24668 );
    not g20061 ( n7723 , n27129 );
    not g20062 ( n11790 , n22442 );
    xnor g20063 ( n23694 , n30895 , n9619 );
    xnor g20064 ( n8454 , n11027 , n24581 );
    not g20065 ( n26855 , n4237 );
    or g20066 ( n681 , n10528 , n19167 );
    not g20067 ( n23050 , n12031 );
    xnor g20068 ( n24607 , n9492 , n6172 );
    not g20069 ( n4817 , n6249 );
    xnor g20070 ( n25580 , n17797 , n29476 );
    not g20071 ( n6448 , n4499 );
    or g20072 ( n31162 , n11841 , n5242 );
    and g20073 ( n7461 , n12973 , n26133 );
    not g20074 ( n3806 , n17761 );
    not g20075 ( n4011 , n3614 );
    nor g20076 ( n6147 , n31326 , n666 );
    not g20077 ( n27258 , n23278 );
    or g20078 ( n2670 , n9417 , n15527 );
    and g20079 ( n16325 , n22965 , n12575 );
    not g20080 ( n5471 , n29764 );
    and g20081 ( n10244 , n4682 , n19824 );
    and g20082 ( n27902 , n14077 , n3551 );
    or g20083 ( n16496 , n5550 , n29546 );
    not g20084 ( n24371 , n8649 );
    or g20085 ( n24154 , n8101 , n11399 );
    and g20086 ( n3137 , n11160 , n26522 );
    or g20087 ( n28881 , n12813 , n26097 );
    and g20088 ( n15280 , n15661 , n23042 );
    and g20089 ( n4814 , n27532 , n2360 );
    xnor g20090 ( n9998 , n5924 , n20486 );
    not g20091 ( n30933 , n10983 );
    xnor g20092 ( n23402 , n21452 , n21918 );
    not g20093 ( n177 , n24324 );
    not g20094 ( n26723 , n18470 );
    not g20095 ( n28103 , n30906 );
    not g20096 ( n18489 , n15827 );
    or g20097 ( n12307 , n22192 , n12780 );
    nor g20098 ( n24680 , n3858 , n12550 );
    xnor g20099 ( n871 , n20911 , n15746 );
    nor g20100 ( n18409 , n7210 , n10842 );
    and g20101 ( n5233 , n28447 , n25175 );
    nor g20102 ( n20750 , n22867 , n24429 );
    and g20103 ( n30730 , n25705 , n18601 );
    xnor g20104 ( n3955 , n13926 , n13899 );
    xnor g20105 ( n15458 , n14489 , n318 );
    or g20106 ( n12583 , n16238 , n13149 );
    and g20107 ( n31423 , n21267 , n7324 );
    not g20108 ( n16056 , n7787 );
    not g20109 ( n1176 , n18470 );
    or g20110 ( n9599 , n15068 , n1340 );
    not g20111 ( n13186 , n20385 );
    or g20112 ( n14448 , n11304 , n3371 );
    nor g20113 ( n3874 , n10927 , n18794 );
    or g20114 ( n6007 , n11065 , n23667 );
    not g20115 ( n6154 , n15397 );
    and g20116 ( n14737 , n3128 , n17351 );
    xnor g20117 ( n21836 , n8422 , n5062 );
    xor g20118 ( n19727 , n14663 , n30195 );
    or g20119 ( n10103 , n31675 , n5524 );
    xnor g20120 ( n22715 , n2345 , n30641 );
    and g20121 ( n26195 , n14229 , n5460 );
    xnor g20122 ( n3411 , n28286 , n28326 );
    not g20123 ( n22778 , n14942 );
    not g20124 ( n17923 , n2019 );
    or g20125 ( n26145 , n4839 , n29813 );
    nor g20126 ( n15324 , n24289 , n3709 );
    and g20127 ( n10354 , n4198 , n16549 );
    not g20128 ( n22745 , n28397 );
    not g20129 ( n5569 , n8791 );
    not g20130 ( n1426 , n10378 );
    nor g20131 ( n8914 , n6195 , n8783 );
    or g20132 ( n24997 , n22760 , n30966 );
    or g20133 ( n14957 , n3345 , n18549 );
    and g20134 ( n24673 , n9351 , n27546 );
    xnor g20135 ( n14858 , n31393 , n4966 );
    and g20136 ( n23427 , n20641 , n26083 );
    and g20137 ( n25750 , n22728 , n1412 );
    not g20138 ( n20106 , n30162 );
    or g20139 ( n13610 , n11999 , n19087 );
    xnor g20140 ( n374 , n5246 , n30651 );
    not g20141 ( n27121 , n5783 );
    not g20142 ( n30467 , n7241 );
    nor g20143 ( n2435 , n31917 , n26577 );
    nor g20144 ( n2394 , n24704 , n29197 );
    or g20145 ( n24295 , n7794 , n18737 );
    not g20146 ( n23927 , n13488 );
    or g20147 ( n15561 , n9358 , n8623 );
    buf g20148 ( n28192 , n12160 );
    not g20149 ( n25265 , n20632 );
    xnor g20150 ( n22971 , n17681 , n19847 );
    xnor g20151 ( n21249 , n16048 , n28901 );
    and g20152 ( n29904 , n7194 , n2688 );
    or g20153 ( n24861 , n22917 , n3080 );
    and g20154 ( n15569 , n30143 , n3424 );
    xnor g20155 ( n28613 , n6161 , n18244 );
    xnor g20156 ( n6474 , n830 , n11462 );
    or g20157 ( n24754 , n9381 , n8767 );
    not g20158 ( n24121 , n18507 );
    xnor g20159 ( n31933 , n17254 , n10676 );
    not g20160 ( n4183 , n28267 );
    not g20161 ( n30516 , n4037 );
    xnor g20162 ( n22368 , n1639 , n30089 );
    and g20163 ( n947 , n17423 , n16693 );
    xnor g20164 ( n12507 , n29438 , n22548 );
    not g20165 ( n4754 , n7163 );
    xnor g20166 ( n20063 , n13624 , n11074 );
    and g20167 ( n17788 , n19354 , n15238 );
    xnor g20168 ( n9966 , n7050 , n28945 );
    not g20169 ( n13865 , n15526 );
    and g20170 ( n7971 , n8070 , n27417 );
    not g20171 ( n8238 , n25695 );
    and g20172 ( n1978 , n178 , n24237 );
    or g20173 ( n25736 , n26598 , n16625 );
    not g20174 ( n7717 , n18829 );
    or g20175 ( n2880 , n17732 , n23940 );
    or g20176 ( n6563 , n14091 , n7901 );
    xnor g20177 ( n5533 , n17656 , n7369 );
    nor g20178 ( n27944 , n8191 , n11979 );
    or g20179 ( n30091 , n5389 , n9304 );
    xnor g20180 ( n8574 , n30499 , n5197 );
    or g20181 ( n25915 , n16268 , n27828 );
    not g20182 ( n11030 , n3540 );
    xnor g20183 ( n7346 , n16129 , n24900 );
    not g20184 ( n16023 , n29836 );
    nor g20185 ( n21957 , n29733 , n21464 );
    or g20186 ( n7924 , n8891 , n22982 );
    and g20187 ( n874 , n8382 , n4279 );
    not g20188 ( n26049 , n19200 );
    xor g20189 ( n7491 , n26577 , n21424 );
    not g20190 ( n2841 , n25389 );
    not g20191 ( n19488 , n8543 );
    and g20192 ( n20945 , n6447 , n4100 );
    xnor g20193 ( n3392 , n17209 , n4213 );
    xnor g20194 ( n3385 , n8048 , n2179 );
    xnor g20195 ( n8811 , n6350 , n22919 );
    nor g20196 ( n12155 , n30529 , n25239 );
    or g20197 ( n20618 , n5146 , n5090 );
    and g20198 ( n748 , n15920 , n5991 );
    or g20199 ( n16118 , n9670 , n21707 );
    not g20200 ( n28410 , n3983 );
    and g20201 ( n7772 , n25652 , n15643 );
    xnor g20202 ( n24691 , n5590 , n24618 );
    xnor g20203 ( n28952 , n12203 , n31186 );
    nor g20204 ( n24911 , n12398 , n27002 );
    xnor g20205 ( n26839 , n11455 , n23650 );
    xnor g20206 ( n1815 , n2961 , n3730 );
    xnor g20207 ( n30957 , n6845 , n3728 );
    not g20208 ( n4174 , n9744 );
    not g20209 ( n4113 , n19717 );
    and g20210 ( n10016 , n7463 , n3104 );
    not g20211 ( n30585 , n645 );
    or g20212 ( n13687 , n31146 , n2538 );
    or g20213 ( n16995 , n18264 , n31325 );
    not g20214 ( n19977 , n26444 );
    nor g20215 ( n23268 , n20118 , n14495 );
    not g20216 ( n11045 , n6211 );
    not g20217 ( n16624 , n3068 );
    and g20218 ( n382 , n19073 , n19715 );
    xnor g20219 ( n5668 , n3819 , n5001 );
    not g20220 ( n11807 , n15733 );
    not g20221 ( n20334 , n9619 );
    not g20222 ( n9505 , n12052 );
    not g20223 ( n28286 , n3596 );
    xnor g20224 ( n22352 , n27014 , n29242 );
    and g20225 ( n6673 , n16169 , n8041 );
    or g20226 ( n13728 , n6249 , n1841 );
    not g20227 ( n10494 , n14656 );
    not g20228 ( n11788 , n2023 );
    nor g20229 ( n29339 , n14555 , n26235 );
    or g20230 ( n11621 , n7435 , n29348 );
    or g20231 ( n706 , n2763 , n4761 );
    not g20232 ( n18302 , n2033 );
    or g20233 ( n19719 , n5116 , n28092 );
    xnor g20234 ( n5011 , n874 , n7824 );
    nor g20235 ( n22752 , n13411 , n3148 );
    or g20236 ( n31925 , n1066 , n8326 );
    nor g20237 ( n15281 , n16132 , n891 );
    and g20238 ( n2492 , n15489 , n17865 );
    not g20239 ( n15397 , n28460 );
    not g20240 ( n820 , n947 );
    not g20241 ( n5327 , n13287 );
    xnor g20242 ( n12518 , n1575 , n8584 );
    not g20243 ( n22300 , n21524 );
    not g20244 ( n22501 , n1559 );
    xnor g20245 ( n27768 , n17149 , n3131 );
    or g20246 ( n23609 , n18552 , n31506 );
    not g20247 ( n24465 , n23559 );
    nor g20248 ( n6146 , n16672 , n265 );
    not g20249 ( n14648 , n7651 );
    or g20250 ( n31569 , n19917 , n1015 );
    and g20251 ( n17098 , n20953 , n22635 );
    not g20252 ( n15110 , n15289 );
    or g20253 ( n29130 , n3670 , n22261 );
    or g20254 ( n18173 , n22234 , n24180 );
    nor g20255 ( n6189 , n26541 , n19100 );
    xnor g20256 ( n31212 , n10826 , n5948 );
    xnor g20257 ( n27327 , n10277 , n19260 );
    or g20258 ( n18341 , n29038 , n16037 );
    xnor g20259 ( n6383 , n6579 , n8388 );
    not g20260 ( n22793 , n14392 );
    or g20261 ( n22772 , n4844 , n10131 );
    nor g20262 ( n15468 , n16088 , n16559 );
    xnor g20263 ( n7833 , n19241 , n13461 );
    or g20264 ( n3376 , n23460 , n30942 );
    xnor g20265 ( n24567 , n15662 , n11708 );
    not g20266 ( n18351 , n18211 );
    or g20267 ( n14797 , n20644 , n13495 );
    xnor g20268 ( n27112 , n12400 , n30669 );
    not g20269 ( n14225 , n8137 );
    not g20270 ( n7860 , n4479 );
    xnor g20271 ( n24557 , n18452 , n22184 );
    not g20272 ( n5242 , n26491 );
    or g20273 ( n13617 , n14925 , n14135 );
    not g20274 ( n25506 , n11789 );
    xnor g20275 ( n24634 , n2535 , n22393 );
    xnor g20276 ( n25152 , n24475 , n19847 );
    or g20277 ( n23929 , n20940 , n22595 );
    xnor g20278 ( n23522 , n12709 , n8617 );
    not g20279 ( n20791 , n6139 );
    not g20280 ( n22951 , n278 );
    not g20281 ( n23626 , n10684 );
    and g20282 ( n17636 , n29749 , n22823 );
    not g20283 ( n7907 , n19494 );
    and g20284 ( n28690 , n24156 , n29250 );
    or g20285 ( n24562 , n1431 , n24231 );
    or g20286 ( n11542 , n7318 , n30380 );
    xnor g20287 ( n21950 , n22995 , n28491 );
    nor g20288 ( n25707 , n21616 , n19283 );
    or g20289 ( n2561 , n26705 , n24444 );
    not g20290 ( n1691 , n30724 );
    xnor g20291 ( n9477 , n23203 , n15977 );
    or g20292 ( n17144 , n17417 , n18260 );
    nor g20293 ( n25933 , n22567 , n24675 );
    xnor g20294 ( n21552 , n2640 , n17305 );
    not g20295 ( n12388 , n1702 );
    and g20296 ( n18240 , n10501 , n27292 );
    or g20297 ( n7867 , n11094 , n1157 );
    or g20298 ( n9425 , n25859 , n19216 );
    nor g20299 ( n18317 , n6874 , n184 );
    not g20300 ( n11676 , n8454 );
    not g20301 ( n3429 , n28545 );
    nor g20302 ( n16538 , n18410 , n9879 );
    and g20303 ( n12671 , n27078 , n20189 );
    xnor g20304 ( n9634 , n18645 , n31773 );
    and g20305 ( n14406 , n23729 , n28823 );
    not g20306 ( n11492 , n20453 );
    xnor g20307 ( n15133 , n9874 , n27278 );
    not g20308 ( n10563 , n3036 );
    or g20309 ( n7300 , n20318 , n25856 );
    not g20310 ( n17898 , n19720 );
    xnor g20311 ( n15779 , n25269 , n25690 );
    or g20312 ( n1958 , n6006 , n20895 );
    xnor g20313 ( n24067 , n26485 , n13043 );
    not g20314 ( n12558 , n30384 );
    xnor g20315 ( n5034 , n29860 , n20342 );
    xnor g20316 ( n22009 , n1832 , n15322 );
    and g20317 ( n26784 , n2157 , n2028 );
    or g20318 ( n22214 , n9902 , n301 );
    or g20319 ( n26081 , n30441 , n29030 );
    and g20320 ( n20416 , n19280 , n8410 );
    not g20321 ( n29546 , n13420 );
    or g20322 ( n11843 , n9239 , n8188 );
    xnor g20323 ( n16043 , n26869 , n11169 );
    or g20324 ( n7826 , n179 , n344 );
    not g20325 ( n1193 , n22057 );
    not g20326 ( n13707 , n9435 );
    and g20327 ( n8231 , n29892 , n10410 );
    not g20328 ( n13152 , n2809 );
    nor g20329 ( n12064 , n26786 , n1032 );
    and g20330 ( n19244 , n10300 , n10646 );
    xor g20331 ( n15663 , n10462 , n15048 );
    not g20332 ( n31636 , n22197 );
    and g20333 ( n321 , n24172 , n11687 );
    or g20334 ( n19180 , n7054 , n23397 );
    not g20335 ( n3266 , n17219 );
    nor g20336 ( n9607 , n30554 , n3711 );
    or g20337 ( n13569 , n14002 , n6065 );
    not g20338 ( n14343 , n28046 );
    or g20339 ( n25410 , n18843 , n18251 );
    nor g20340 ( n1423 , n31108 , n6072 );
    not g20341 ( n12696 , n19456 );
    not g20342 ( n4757 , n11760 );
    not g20343 ( n16135 , n9239 );
    not g20344 ( n2719 , n31470 );
    or g20345 ( n2131 , n24023 , n7277 );
    not g20346 ( n20318 , n21597 );
    or g20347 ( n19278 , n20325 , n8725 );
    and g20348 ( n23039 , n27212 , n15581 );
    not g20349 ( n21606 , n6172 );
    and g20350 ( n21415 , n127 , n25086 );
    not g20351 ( n3506 , n20312 );
    and g20352 ( n24017 , n22404 , n12499 );
    xnor g20353 ( n24356 , n4182 , n641 );
    and g20354 ( n21029 , n10820 , n9580 );
    not g20355 ( n27747 , n17077 );
    nor g20356 ( n15096 , n22294 , n12084 );
    xnor g20357 ( n1574 , n21992 , n22865 );
    nor g20358 ( n29292 , n19208 , n16117 );
    not g20359 ( n29568 , n20495 );
    or g20360 ( n28949 , n23229 , n7610 );
    or g20361 ( n31238 , n8077 , n23330 );
    not g20362 ( n6125 , n9653 );
    not g20363 ( n21993 , n13171 );
    nor g20364 ( n20880 , n6397 , n3015 );
    not g20365 ( n7319 , n9609 );
    xnor g20366 ( n10262 , n25362 , n953 );
    not g20367 ( n2734 , n26894 );
    xnor g20368 ( n2010 , n13381 , n22689 );
    or g20369 ( n10752 , n28023 , n15031 );
    nor g20370 ( n13025 , n14373 , n11755 );
    not g20371 ( n18331 , n25581 );
    or g20372 ( n4518 , n7522 , n12286 );
    xnor g20373 ( n11390 , n25318 , n1241 );
    not g20374 ( n23818 , n16033 );
    nor g20375 ( n16445 , n27580 , n9438 );
    xor g20376 ( n25273 , n9965 , n24167 );
    nor g20377 ( n22012 , n27020 , n10569 );
    not g20378 ( n1806 , n1569 );
    or g20379 ( n12357 , n26383 , n12029 );
    or g20380 ( n5482 , n7883 , n28538 );
    not g20381 ( n13348 , n13591 );
    and g20382 ( n1385 , n13118 , n10891 );
    xnor g20383 ( n650 , n28856 , n3268 );
    not g20384 ( n11491 , n12610 );
    and g20385 ( n3857 , n15801 , n11831 );
    xnor g20386 ( n25308 , n14802 , n28063 );
    not g20387 ( n26033 , n20504 );
    xnor g20388 ( n15278 , n16133 , n18676 );
    not g20389 ( n6278 , n5086 );
    not g20390 ( n12405 , n3117 );
    and g20391 ( n8176 , n24025 , n19543 );
    not g20392 ( n14233 , n22747 );
    xnor g20393 ( n15751 , n11116 , n11692 );
    xor g20394 ( n2960 , n24910 , n2544 );
    and g20395 ( n6124 , n17799 , n30844 );
    not g20396 ( n27911 , n8967 );
    and g20397 ( n12039 , n25256 , n30138 );
    and g20398 ( n30212 , n20294 , n10487 );
    buf g20399 ( n30813 , n16250 );
    xor g20400 ( n31945 , n16792 , n18392 );
    or g20401 ( n11444 , n23047 , n1351 );
    nor g20402 ( n16366 , n15719 , n12934 );
    nor g20403 ( n23141 , n26404 , n13788 );
    not g20404 ( n26905 , n975 );
    and g20405 ( n8679 , n11240 , n7045 );
    nor g20406 ( n24408 , n9948 , n16238 );
    not g20407 ( n17547 , n15195 );
    xnor g20408 ( n3086 , n7205 , n3312 );
    and g20409 ( n24150 , n12667 , n7578 );
    xnor g20410 ( n27230 , n15152 , n12867 );
    not g20411 ( n285 , n13983 );
    nor g20412 ( n30377 , n11850 , n24574 );
    xnor g20413 ( n23288 , n821 , n5484 );
    and g20414 ( n16984 , n15332 , n4195 );
    xor g20415 ( n6840 , n10091 , n14954 );
    xnor g20416 ( n19517 , n4695 , n739 );
    and g20417 ( n5835 , n2659 , n16919 );
    not g20418 ( n8735 , n9334 );
    xnor g20419 ( n5680 , n16459 , n18282 );
    not g20420 ( n6449 , n2431 );
    xnor g20421 ( n20726 , n25418 , n27206 );
    not g20422 ( n29095 , n29132 );
    not g20423 ( n31713 , n3587 );
    xnor g20424 ( n7648 , n20202 , n17427 );
    or g20425 ( n7554 , n17149 , n4701 );
    or g20426 ( n3944 , n1980 , n14861 );
    not g20427 ( n30724 , n2550 );
    not g20428 ( n6149 , n2923 );
    xnor g20429 ( n471 , n22153 , n18534 );
    or g20430 ( n7185 , n30970 , n8598 );
    not g20431 ( n13665 , n16031 );
    nor g20432 ( n16005 , n7218 , n1870 );
    not g20433 ( n24833 , n11635 );
    not g20434 ( n10845 , n10019 );
    or g20435 ( n16818 , n2110 , n5292 );
    xor g20436 ( n21612 , n11517 , n3277 );
    not g20437 ( n25904 , n29569 );
    not g20438 ( n31847 , n26114 );
    or g20439 ( n25471 , n29183 , n23867 );
    not g20440 ( n25336 , n13122 );
    not g20441 ( n21636 , n27613 );
    not g20442 ( n25616 , n28748 );
    nor g20443 ( n15784 , n23897 , n26327 );
    or g20444 ( n8312 , n15884 , n13741 );
    xnor g20445 ( n1844 , n2279 , n15174 );
    xnor g20446 ( n17452 , n10368 , n1876 );
    xnor g20447 ( n488 , n20839 , n3710 );
    or g20448 ( n27450 , n25443 , n30879 );
    or g20449 ( n25642 , n22047 , n23112 );
    and g20450 ( n5081 , n14756 , n27097 );
    not g20451 ( n19907 , n12922 );
    nor g20452 ( n30494 , n12874 , n9094 );
    and g20453 ( n13915 , n11001 , n22700 );
    or g20454 ( n24740 , n5251 , n8189 );
    not g20455 ( n1334 , n26220 );
    xnor g20456 ( n359 , n22615 , n6380 );
    and g20457 ( n760 , n4745 , n3203 );
    not g20458 ( n26583 , n30758 );
    or g20459 ( n20965 , n27974 , n24232 );
    not g20460 ( n20530 , n12797 );
    nor g20461 ( n21329 , n7854 , n23189 );
    xnor g20462 ( n15454 , n27087 , n26957 );
    xnor g20463 ( n13708 , n27475 , n13526 );
    not g20464 ( n2378 , n4604 );
    and g20465 ( n29934 , n7225 , n27951 );
    xnor g20466 ( n328 , n13499 , n18749 );
    not g20467 ( n9242 , n11339 );
    nor g20468 ( n16349 , n17291 , n16061 );
    not g20469 ( n11017 , n19765 );
    xnor g20470 ( n19841 , n20942 , n854 );
    and g20471 ( n2771 , n9972 , n9408 );
    xnor g20472 ( n14794 , n17413 , n25261 );
    nor g20473 ( n413 , n2925 , n1095 );
    and g20474 ( n31879 , n19417 , n2891 );
    xnor g20475 ( n29159 , n7902 , n5293 );
    and g20476 ( n2295 , n1287 , n28079 );
    and g20477 ( n2015 , n19145 , n16877 );
    nor g20478 ( n19835 , n7692 , n24487 );
    xnor g20479 ( n22281 , n17391 , n13618 );
    nor g20480 ( n26531 , n17499 , n30036 );
    not g20481 ( n10838 , n12409 );
    or g20482 ( n8481 , n31942 , n10703 );
    nor g20483 ( n14291 , n21141 , n23127 );
    or g20484 ( n14948 , n8713 , n24068 );
    and g20485 ( n14570 , n12909 , n17975 );
    xnor g20486 ( n12261 , n15807 , n23043 );
    not g20487 ( n2225 , n318 );
    or g20488 ( n6025 , n30831 , n5451 );
    xnor g20489 ( n16672 , n22754 , n17227 );
    and g20490 ( n10967 , n10020 , n2118 );
    not g20491 ( n15584 , n7314 );
    not g20492 ( n7362 , n4414 );
    xnor g20493 ( n20351 , n10332 , n21963 );
    or g20494 ( n6699 , n14791 , n15415 );
    not g20495 ( n17029 , n10134 );
    and g20496 ( n28414 , n16519 , n16646 );
    and g20497 ( n482 , n4578 , n819 );
    xnor g20498 ( n25500 , n4278 , n6349 );
    xnor g20499 ( n22664 , n7306 , n477 );
    and g20500 ( n22494 , n26079 , n8519 );
    nor g20501 ( n2774 , n15917 , n22256 );
    or g20502 ( n403 , n22423 , n27591 );
    xnor g20503 ( n31473 , n11717 , n21685 );
    or g20504 ( n5238 , n20907 , n20143 );
    nor g20505 ( n27123 , n12112 , n10674 );
    not g20506 ( n24116 , n5986 );
    xnor g20507 ( n29682 , n21182 , n16685 );
    xnor g20508 ( n2494 , n12436 , n15223 );
    and g20509 ( n11033 , n19126 , n29959 );
    not g20510 ( n21242 , n1567 );
    not g20511 ( n20968 , n2950 );
    and g20512 ( n24231 , n23783 , n10678 );
    xnor g20513 ( n16417 , n25527 , n19132 );
    xnor g20514 ( n27528 , n15817 , n28909 );
    and g20515 ( n23447 , n5184 , n24342 );
    not g20516 ( n29781 , n17044 );
    xnor g20517 ( n16310 , n8208 , n12777 );
    xnor g20518 ( n18134 , n22588 , n1629 );
    and g20519 ( n23070 , n21012 , n28768 );
    not g20520 ( n19598 , n30271 );
    xnor g20521 ( n6399 , n15518 , n4917 );
    or g20522 ( n9893 , n12207 , n8897 );
    not g20523 ( n15289 , n10904 );
    and g20524 ( n20985 , n29577 , n14146 );
    not g20525 ( n13838 , n24546 );
    not g20526 ( n25715 , n25426 );
    not g20527 ( n12377 , n25108 );
    or g20528 ( n8519 , n8249 , n29658 );
    or g20529 ( n7486 , n19508 , n25162 );
    xnor g20530 ( n10130 , n2815 , n2021 );
    nor g20531 ( n19074 , n22139 , n25543 );
    not g20532 ( n1872 , n4308 );
    and g20533 ( n4738 , n30760 , n1533 );
    and g20534 ( n1099 , n21219 , n26645 );
    not g20535 ( n28173 , n5951 );
    nor g20536 ( n2721 , n2221 , n21549 );
    and g20537 ( n261 , n3556 , n19827 );
    or g20538 ( n23221 , n11103 , n23241 );
    not g20539 ( n24171 , n25757 );
    not g20540 ( n23258 , n10451 );
    xnor g20541 ( n29589 , n30812 , n5638 );
    or g20542 ( n2647 , n21536 , n14778 );
    and g20543 ( n24099 , n7373 , n13377 );
    or g20544 ( n25566 , n28400 , n10516 );
    or g20545 ( n1326 , n9942 , n5468 );
    not g20546 ( n8363 , n6349 );
    xnor g20547 ( n13043 , n8257 , n4697 );
    xnor g20548 ( n1063 , n8412 , n14615 );
    xor g20549 ( n5131 , n5735 , n14667 );
    not g20550 ( n30352 , n8421 );
    nor g20551 ( n994 , n12349 , n8363 );
    and g20552 ( n13087 , n31101 , n5407 );
    not g20553 ( n25563 , n14303 );
    or g20554 ( n88 , n18283 , n25227 );
    or g20555 ( n19417 , n18225 , n16542 );
    or g20556 ( n21526 , n18960 , n27729 );
    nor g20557 ( n20974 , n11421 , n13357 );
    nor g20558 ( n29097 , n7253 , n11823 );
    not g20559 ( n10888 , n22262 );
    xnor g20560 ( n10699 , n1092 , n31021 );
    and g20561 ( n21740 , n30492 , n5158 );
    or g20562 ( n14581 , n20278 , n17299 );
    or g20563 ( n3697 , n7012 , n29473 );
    xnor g20564 ( n15422 , n11841 , n26963 );
    xnor g20565 ( n19385 , n23115 , n16075 );
    and g20566 ( n4763 , n31459 , n31852 );
    and g20567 ( n8671 , n24159 , n4838 );
    or g20568 ( n9068 , n19426 , n29690 );
    or g20569 ( n10754 , n8208 , n17663 );
    xnor g20570 ( n3248 , n23762 , n6137 );
    not g20571 ( n16094 , n8282 );
    nor g20572 ( n1609 , n28951 , n15829 );
    not g20573 ( n24002 , n17302 );
    not g20574 ( n26948 , n18042 );
    xnor g20575 ( n27150 , n28108 , n4650 );
    xnor g20576 ( n24879 , n6825 , n290 );
    and g20577 ( n7585 , n26497 , n4835 );
    xnor g20578 ( n1960 , n1865 , n1331 );
    nor g20579 ( n14352 , n2311 , n30867 );
    xnor g20580 ( n18905 , n16955 , n26292 );
    xnor g20581 ( n13829 , n7516 , n7518 );
    xnor g20582 ( n11829 , n10427 , n14688 );
    or g20583 ( n10824 , n10166 , n30460 );
    xnor g20584 ( n22007 , n12015 , n19979 );
    xnor g20585 ( n13239 , n12344 , n21540 );
    xnor g20586 ( n28774 , n10530 , n5183 );
    and g20587 ( n22051 , n20674 , n1828 );
    not g20588 ( n14473 , n7296 );
    and g20589 ( n6990 , n1503 , n22102 );
    not g20590 ( n10634 , n16238 );
    buf g20591 ( n26264 , n21717 );
    xnor g20592 ( n13705 , n13576 , n3596 );
    xnor g20593 ( n3844 , n23026 , n11913 );
    xnor g20594 ( n12392 , n19403 , n13940 );
    or g20595 ( n7519 , n23047 , n26748 );
    or g20596 ( n18324 , n27801 , n10284 );
    xnor g20597 ( n21455 , n2114 , n31445 );
    not g20598 ( n23550 , n3169 );
    or g20599 ( n25656 , n9386 , n24771 );
    or g20600 ( n20182 , n13572 , n15373 );
    not g20601 ( n4072 , n30534 );
    nor g20602 ( n22609 , n22163 , n1172 );
    and g20603 ( n19559 , n6402 , n9588 );
    or g20604 ( n3201 , n18968 , n14856 );
    xnor g20605 ( n3580 , n25027 , n27089 );
    not g20606 ( n12230 , n5443 );
    not g20607 ( n22545 , n10179 );
    nor g20608 ( n1561 , n10413 , n30689 );
    xnor g20609 ( n1917 , n11159 , n7144 );
    and g20610 ( n16616 , n10022 , n13459 );
    and g20611 ( n4286 , n8633 , n12391 );
    xnor g20612 ( n5100 , n30410 , n15802 );
    xnor g20613 ( n30850 , n12398 , n27002 );
    and g20614 ( n12644 , n27915 , n3035 );
    or g20615 ( n14453 , n8668 , n13937 );
    or g20616 ( n24117 , n697 , n7421 );
    and g20617 ( n5928 , n28200 , n6332 );
    and g20618 ( n31628 , n10618 , n30493 );
    xnor g20619 ( n1921 , n61 , n1172 );
    not g20620 ( n2443 , n6226 );
    not g20621 ( n30290 , n11462 );
    and g20622 ( n21396 , n16339 , n6414 );
    xnor g20623 ( n3396 , n18026 , n18907 );
    or g20624 ( n19898 , n319 , n26581 );
    or g20625 ( n17666 , n29090 , n20799 );
    not g20626 ( n22242 , n19770 );
    xnor g20627 ( n25539 , n5427 , n22601 );
    not g20628 ( n8443 , n22731 );
    not g20629 ( n9185 , n28292 );
    and g20630 ( n27397 , n25475 , n31987 );
    xnor g20631 ( n17230 , n28570 , n19780 );
    or g20632 ( n21858 , n28441 , n25254 );
    nor g20633 ( n25264 , n23360 , n6098 );
    xnor g20634 ( n14816 , n11825 , n1276 );
    nor g20635 ( n9483 , n4213 , n3184 );
    xnor g20636 ( n22471 , n5388 , n10327 );
    xnor g20637 ( n1500 , n30358 , n22925 );
    xnor g20638 ( n27696 , n21243 , n7632 );
    xnor g20639 ( n28155 , n23040 , n29090 );
    or g20640 ( n1578 , n16873 , n20181 );
    not g20641 ( n30732 , n17132 );
    not g20642 ( n15214 , n18203 );
    xnor g20643 ( n14979 , n18498 , n21279 );
    nor g20644 ( n25639 , n3080 , n27605 );
    or g20645 ( n14060 , n1302 , n21443 );
    or g20646 ( n25652 , n17106 , n30944 );
    nor g20647 ( n10746 , n10014 , n21537 );
    or g20648 ( n7294 , n2756 , n6670 );
    xnor g20649 ( n2235 , n16142 , n31305 );
    and g20650 ( n13830 , n1185 , n28343 );
    xnor g20651 ( n13004 , n4989 , n9077 );
    nor g20652 ( n26023 , n16345 , n14766 );
    xnor g20653 ( n8130 , n31070 , n28828 );
    and g20654 ( n24818 , n25126 , n18294 );
    xnor g20655 ( n18977 , n3148 , n24943 );
    and g20656 ( n8032 , n14749 , n4558 );
    or g20657 ( n22312 , n3648 , n2922 );
    and g20658 ( n6670 , n23009 , n2945 );
    nor g20659 ( n16282 , n30449 , n16828 );
    not g20660 ( n19521 , n16264 );
    and g20661 ( n25523 , n5225 , n2254 );
    and g20662 ( n13422 , n25216 , n9990 );
    or g20663 ( n8243 , n395 , n25755 );
    or g20664 ( n1996 , n20997 , n11511 );
    not g20665 ( n13046 , n22551 );
    xnor g20666 ( n9961 , n17603 , n16225 );
    xnor g20667 ( n18769 , n25982 , n27805 );
    not g20668 ( n7940 , n687 );
    not g20669 ( n996 , n27969 );
    not g20670 ( n2879 , n21771 );
    not g20671 ( n9616 , n18234 );
    not g20672 ( n9345 , n27453 );
    not g20673 ( n2130 , n13664 );
    or g20674 ( n25301 , n16626 , n15602 );
    or g20675 ( n7984 , n15137 , n18122 );
    or g20676 ( n7631 , n26049 , n16578 );
    or g20677 ( n5738 , n5751 , n27314 );
    xnor g20678 ( n24167 , n30094 , n6745 );
    xnor g20679 ( n3229 , n4901 , n8133 );
    nor g20680 ( n8061 , n7981 , n3702 );
    nor g20681 ( n27398 , n27355 , n25646 );
    xor g20682 ( n17195 , n13508 , n20815 );
    or g20683 ( n30332 , n26709 , n18308 );
    and g20684 ( n17637 , n1855 , n4870 );
    nor g20685 ( n12753 , n10045 , n26233 );
    xnor g20686 ( n29106 , n24190 , n1982 );
    or g20687 ( n14935 , n25529 , n21415 );
    or g20688 ( n29894 , n19773 , n9955 );
    xnor g20689 ( n29261 , n25713 , n28745 );
    or g20690 ( n7868 , n238 , n13752 );
    or g20691 ( n12206 , n320 , n29036 );
    and g20692 ( n20462 , n25347 , n20155 );
    not g20693 ( n24758 , n13990 );
    not g20694 ( n10792 , n28243 );
    xnor g20695 ( n13215 , n17297 , n17196 );
    and g20696 ( n31803 , n17576 , n28895 );
    xnor g20697 ( n20933 , n28102 , n7692 );
    and g20698 ( n19039 , n29220 , n1729 );
    and g20699 ( n5774 , n5210 , n12599 );
    and g20700 ( n24959 , n22923 , n1992 );
    not g20701 ( n26217 , n24980 );
    nor g20702 ( n12665 , n29615 , n10259 );
    xnor g20703 ( n21107 , n3672 , n17174 );
    not g20704 ( n14846 , n21918 );
    not g20705 ( n8742 , n1284 );
    not g20706 ( n25280 , n24582 );
    and g20707 ( n25304 , n17420 , n8106 );
    or g20708 ( n28859 , n8241 , n562 );
    or g20709 ( n19129 , n4173 , n24479 );
    and g20710 ( n30210 , n29794 , n17413 );
    and g20711 ( n14219 , n26395 , n23884 );
    not g20712 ( n27863 , n15532 );
    not g20713 ( n17289 , n8867 );
    and g20714 ( n2065 , n29042 , n21161 );
    not g20715 ( n29145 , n18598 );
    xnor g20716 ( n31413 , n24953 , n31940 );
    not g20717 ( n7330 , n11071 );
    xor g20718 ( n24482 , n20017 , n14563 );
    not g20719 ( n4532 , n28169 );
    xnor g20720 ( n4175 , n25782 , n15751 );
    xnor g20721 ( n29732 , n15885 , n27970 );
    not g20722 ( n13658 , n28923 );
    xnor g20723 ( n17575 , n19050 , n13601 );
    or g20724 ( n13251 , n30023 , n91 );
    not g20725 ( n7623 , n25670 );
    nor g20726 ( n20250 , n7210 , n13378 );
    or g20727 ( n30417 , n13720 , n24959 );
    not g20728 ( n2218 , n8195 );
    and g20729 ( n2344 , n19932 , n13435 );
    or g20730 ( n16051 , n20672 , n8409 );
    not g20731 ( n31812 , n7465 );
    not g20732 ( n13174 , n13005 );
    or g20733 ( n18818 , n24730 , n22417 );
    not g20734 ( n6207 , n13539 );
    and g20735 ( n9749 , n6891 , n4309 );
    not g20736 ( n18367 , n28666 );
    or g20737 ( n24810 , n4150 , n6562 );
    and g20738 ( n14750 , n26011 , n3693 );
    and g20739 ( n17555 , n1387 , n22918 );
    or g20740 ( n11464 , n19538 , n31626 );
    or g20741 ( n597 , n23283 , n16057 );
    xnor g20742 ( n17378 , n13320 , n31618 );
    or g20743 ( n7985 , n9267 , n6478 );
    not g20744 ( n23724 , n17491 );
    and g20745 ( n24273 , n12110 , n4985 );
    not g20746 ( n10864 , n1378 );
    or g20747 ( n6790 , n9225 , n14296 );
    or g20748 ( n8492 , n7620 , n20831 );
    or g20749 ( n6764 , n30387 , n23369 );
    or g20750 ( n4293 , n11060 , n31479 );
    or g20751 ( n30652 , n24019 , n26557 );
    or g20752 ( n26802 , n25760 , n3268 );
    xnor g20753 ( n1165 , n18452 , n26306 );
    and g20754 ( n20528 , n31581 , n2941 );
    not g20755 ( n12193 , n4535 );
    nor g20756 ( n18408 , n5382 , n26619 );
    nor g20757 ( n21083 , n7315 , n29897 );
    nor g20758 ( n12658 , n31885 , n14694 );
    and g20759 ( n14605 , n12809 , n24294 );
    xnor g20760 ( n3446 , n13787 , n15325 );
    not g20761 ( n8626 , n21305 );
    xnor g20762 ( n11722 , n2426 , n14930 );
    or g20763 ( n11515 , n26485 , n24294 );
    and g20764 ( n27268 , n9823 , n10919 );
    and g20765 ( n11578 , n16395 , n26448 );
    not g20766 ( n9943 , n30948 );
    xnor g20767 ( n22590 , n23416 , n22139 );
    or g20768 ( n14888 , n13996 , n450 );
    and g20769 ( n1929 , n16127 , n27159 );
    not g20770 ( n14563 , n9825 );
    xnor g20771 ( n14230 , n10613 , n18639 );
    or g20772 ( n20806 , n26092 , n29094 );
    or g20773 ( n30868 , n21019 , n22344 );
    not g20774 ( n27784 , n14557 );
    or g20775 ( n23894 , n1965 , n21495 );
    and g20776 ( n7680 , n27463 , n19338 );
    not g20777 ( n6912 , n1615 );
    not g20778 ( n30553 , n14121 );
    not g20779 ( n6170 , n27500 );
    xnor g20780 ( n19146 , n25317 , n16813 );
    or g20781 ( n30973 , n19211 , n30927 );
    or g20782 ( n5423 , n3510 , n26586 );
    not g20783 ( n26337 , n19221 );
    xnor g20784 ( n19124 , n13149 , n16238 );
    or g20785 ( n25322 , n14112 , n6867 );
    or g20786 ( n29658 , n31 , n20109 );
    xnor g20787 ( n5026 , n9383 , n21422 );
    and g20788 ( n21387 , n5501 , n20226 );
    nor g20789 ( n29156 , n22324 , n16393 );
    not g20790 ( n1485 , n18336 );
    or g20791 ( n31860 , n14773 , n6418 );
    and g20792 ( n20381 , n23177 , n32007 );
    not g20793 ( n4588 , n8439 );
    and g20794 ( n15889 , n11241 , n23842 );
    xnor g20795 ( n4270 , n26717 , n5580 );
    not g20796 ( n13221 , n15320 );
    xnor g20797 ( n31662 , n3322 , n5924 );
    xnor g20798 ( n19596 , n16532 , n1448 );
    and g20799 ( n16117 , n19638 , n11126 );
    not g20800 ( n19693 , n22867 );
    and g20801 ( n24645 , n11744 , n5206 );
    xnor g20802 ( n26534 , n1548 , n8673 );
    nor g20803 ( n21805 , n3192 , n22906 );
    xnor g20804 ( n20845 , n3973 , n22451 );
    xnor g20805 ( n17692 , n12426 , n12143 );
    xnor g20806 ( n9751 , n18075 , n6852 );
    not g20807 ( n24271 , n13697 );
    nor g20808 ( n7054 , n7974 , n953 );
    or g20809 ( n28792 , n21400 , n23636 );
    not g20810 ( n6209 , n31551 );
    not g20811 ( n2022 , n25524 );
    and g20812 ( n27617 , n4364 , n14501 );
    not g20813 ( n23840 , n4412 );
    xnor g20814 ( n24115 , n8791 , n1113 );
    not g20815 ( n15044 , n7745 );
    xnor g20816 ( n28510 , n17469 , n27394 );
    or g20817 ( n22308 , n9930 , n30483 );
    xnor g20818 ( n10703 , n8212 , n20437 );
    nor g20819 ( n26488 , n14670 , n7465 );
    not g20820 ( n13378 , n9655 );
    xnor g20821 ( n29540 , n6348 , n27937 );
    xnor g20822 ( n6734 , n17507 , n1198 );
    and g20823 ( n22676 , n2452 , n1310 );
    not g20824 ( n7732 , n30707 );
    nor g20825 ( n16944 , n17469 , n27394 );
    xnor g20826 ( n19738 , n8946 , n1528 );
    not g20827 ( n9530 , n9531 );
    or g20828 ( n15200 , n30132 , n24492 );
    xnor g20829 ( n3139 , n18044 , n5536 );
    and g20830 ( n29778 , n27611 , n6011 );
    nor g20831 ( n12632 , n27829 , n13972 );
    not g20832 ( n28509 , n30556 );
    xnor g20833 ( n5672 , n28667 , n26346 );
    not g20834 ( n30160 , n5405 );
    or g20835 ( n29247 , n3693 , n26011 );
    or g20836 ( n19789 , n19586 , n29155 );
    xnor g20837 ( n85 , n28539 , n6369 );
    nor g20838 ( n9154 , n29437 , n24687 );
    and g20839 ( n15279 , n2783 , n22884 );
    not g20840 ( n31652 , n32024 );
    xor g20841 ( n13225 , n15020 , n3297 );
    or g20842 ( n26642 , n18616 , n21042 );
    or g20843 ( n20239 , n10374 , n1522 );
    or g20844 ( n10670 , n24377 , n28113 );
    not g20845 ( n6311 , n4092 );
    xnor g20846 ( n547 , n20794 , n14079 );
    xnor g20847 ( n10171 , n12137 , n30659 );
    nor g20848 ( n12954 , n29649 , n26467 );
    not g20849 ( n12184 , n5912 );
    or g20850 ( n6266 , n26318 , n656 );
    or g20851 ( n21431 , n10032 , n7017 );
    not g20852 ( n18058 , n24573 );
    and g20853 ( n26209 , n15513 , n29634 );
    and g20854 ( n21698 , n19020 , n3525 );
    xnor g20855 ( n1630 , n29745 , n10676 );
    and g20856 ( n10286 , n14266 , n7046 );
    not g20857 ( n12522 , n10614 );
    and g20858 ( n24125 , n20003 , n27727 );
    xnor g20859 ( n1118 , n3214 , n22675 );
    and g20860 ( n6828 , n15692 , n8080 );
    xnor g20861 ( n25740 , n28398 , n454 );
    xnor g20862 ( n115 , n10707 , n624 );
    not g20863 ( n20252 , n24086 );
    not g20864 ( n17746 , n27233 );
    not g20865 ( n17265 , n16457 );
    and g20866 ( n2947 , n22249 , n13452 );
    not g20867 ( n2334 , n15190 );
    xnor g20868 ( n7551 , n9147 , n28227 );
    or g20869 ( n30827 , n21311 , n920 );
    or g20870 ( n12375 , n7376 , n74 );
    not g20871 ( n4488 , n10905 );
    or g20872 ( n20648 , n9591 , n26413 );
    not g20873 ( n3361 , n7225 );
    or g20874 ( n9214 , n6067 , n23702 );
    and g20875 ( n27577 , n25643 , n4847 );
    xnor g20876 ( n13690 , n17742 , n84 );
    xnor g20877 ( n31839 , n8801 , n28836 );
    xor g20878 ( n9135 , n6820 , n8955 );
    or g20879 ( n4281 , n22030 , n4455 );
    xnor g20880 ( n11967 , n27773 , n4913 );
    xnor g20881 ( n19138 , n14967 , n24304 );
    xnor g20882 ( n31618 , n16724 , n13338 );
    and g20883 ( n31452 , n8725 , n31415 );
    xnor g20884 ( n17126 , n9331 , n4510 );
    or g20885 ( n25356 , n30690 , n23484 );
    xnor g20886 ( n19331 , n5849 , n22534 );
    xor g20887 ( n2563 , n2476 , n28603 );
    not g20888 ( n1748 , n12028 );
    not g20889 ( n21450 , n22996 );
    not g20890 ( n14485 , n12628 );
    and g20891 ( n23289 , n19691 , n23888 );
    or g20892 ( n9392 , n10139 , n6346 );
    or g20893 ( n25100 , n6936 , n21932 );
    xnor g20894 ( n25954 , n22775 , n11169 );
    not g20895 ( n24152 , n14388 );
    xnor g20896 ( n11005 , n11469 , n24291 );
    not g20897 ( n12710 , n27204 );
    or g20898 ( n20404 , n14875 , n28208 );
    xnor g20899 ( n875 , n4549 , n5793 );
    and g20900 ( n1765 , n19865 , n27569 );
    not g20901 ( n8173 , n25755 );
    or g20902 ( n24862 , n465 , n17926 );
    not g20903 ( n5018 , n16855 );
    xor g20904 ( n15692 , n11071 , n21220 );
    or g20905 ( n19064 , n9715 , n11652 );
    nor g20906 ( n2338 , n13888 , n20859 );
    not g20907 ( n19456 , n2936 );
    not g20908 ( n31013 , n10962 );
    or g20909 ( n30985 , n12428 , n7127 );
    xnor g20910 ( n5493 , n12718 , n26534 );
    or g20911 ( n342 , n12 , n19849 );
    not g20912 ( n6956 , n6658 );
    not g20913 ( n25220 , n12527 );
    nor g20914 ( n6864 , n16947 , n19291 );
    and g20915 ( n21278 , n7061 , n19530 );
    or g20916 ( n25651 , n26712 , n26898 );
    not g20917 ( n29901 , n22096 );
    or g20918 ( n12129 , n29688 , n9349 );
    nor g20919 ( n7500 , n13271 , n27184 );
    not g20920 ( n24728 , n7580 );
    not g20921 ( n6796 , n4840 );
    nor g20922 ( n30818 , n28824 , n24354 );
    or g20923 ( n16754 , n19308 , n24269 );
    not g20924 ( n12890 , n22882 );
    not g20925 ( n3770 , n3491 );
    and g20926 ( n4740 , n21998 , n11933 );
    or g20927 ( n25097 , n30201 , n18166 );
    and g20928 ( n9022 , n31045 , n31871 );
    or g20929 ( n4099 , n25649 , n24520 );
    xnor g20930 ( n3199 , n9716 , n31627 );
    or g20931 ( n3809 , n21292 , n26117 );
    or g20932 ( n24330 , n23115 , n22352 );
    xnor g20933 ( n27643 , n26946 , n28318 );
    not g20934 ( n29003 , n1710 );
    or g20935 ( n9232 , n3680 , n29707 );
    not g20936 ( n18679 , n1931 );
    xnor g20937 ( n27981 , n21059 , n29207 );
    xnor g20938 ( n19346 , n16112 , n27538 );
    or g20939 ( n360 , n31525 , n750 );
    nor g20940 ( n31553 , n590 , n31551 );
    not g20941 ( n1633 , n6236 );
    nor g20942 ( n1370 , n30189 , n5834 );
    not g20943 ( n13436 , n9373 );
    not g20944 ( n1728 , n20428 );
    and g20945 ( n3386 , n20779 , n14091 );
    xnor g20946 ( n1794 , n29312 , n30577 );
    xnor g20947 ( n15878 , n8556 , n298 );
    nor g20948 ( n5811 , n15436 , n12066 );
    and g20949 ( n1536 , n9492 , n21606 );
    not g20950 ( n23861 , n25970 );
    xnor g20951 ( n28359 , n4068 , n31815 );
    xnor g20952 ( n16442 , n183 , n16477 );
    not g20953 ( n31807 , n22170 );
    or g20954 ( n11011 , n10206 , n17282 );
    xnor g20955 ( n2638 , n15498 , n27178 );
    not g20956 ( n13084 , n18048 );
    xnor g20957 ( n11242 , n9627 , n23137 );
    not g20958 ( n19325 , n20607 );
    not g20959 ( n12191 , n15236 );
    or g20960 ( n22334 , n20975 , n10869 );
    or g20961 ( n27165 , n28985 , n17569 );
    and g20962 ( n14986 , n30511 , n20197 );
    not g20963 ( n30189 , n4278 );
    not g20964 ( n11954 , n12074 );
    not g20965 ( n17866 , n29945 );
    not g20966 ( n188 , n21556 );
    xnor g20967 ( n4784 , n3875 , n1278 );
    xnor g20968 ( n27467 , n19253 , n31665 );
    and g20969 ( n10324 , n25656 , n24252 );
    and g20970 ( n13477 , n24559 , n12824 );
    and g20971 ( n11254 , n17323 , n759 );
    xnor g20972 ( n2746 , n5453 , n6438 );
    nor g20973 ( n6683 , n4427 , n7642 );
    or g20974 ( n23958 , n18868 , n30791 );
    not g20975 ( n19512 , n10266 );
    xnor g20976 ( n20549 , n12712 , n18380 );
    xnor g20977 ( n17649 , n7898 , n20278 );
    not g20978 ( n18421 , n7725 );
    xnor g20979 ( n13142 , n17405 , n8030 );
    or g20980 ( n31311 , n15238 , n19354 );
    or g20981 ( n11825 , n11108 , n14038 );
    or g20982 ( n18039 , n19702 , n11555 );
    or g20983 ( n22328 , n13793 , n21992 );
    xnor g20984 ( n5203 , n7587 , n17798 );
    and g20985 ( n21509 , n9637 , n5437 );
    xnor g20986 ( n12438 , n10000 , n19882 );
    xnor g20987 ( n2621 , n14196 , n1819 );
    or g20988 ( n24314 , n27623 , n16158 );
    nor g20989 ( n3296 , n13701 , n16810 );
    not g20990 ( n16316 , n19198 );
    buf g20991 ( n3034 , n23100 );
    or g20992 ( n11061 , n17036 , n5596 );
    or g20993 ( n26875 , n8496 , n25724 );
    nor g20994 ( n19941 , n13145 , n24173 );
    nor g20995 ( n10270 , n891 , n12342 );
    and g20996 ( n18863 , n551 , n11866 );
    or g20997 ( n20448 , n9664 , n26303 );
    nor g20998 ( n11535 , n21646 , n8667 );
    xnor g20999 ( n15991 , n19967 , n31643 );
    and g21000 ( n24729 , n14973 , n17560 );
    xnor g21001 ( n24938 , n18384 , n12273 );
    not g21002 ( n14895 , n9399 );
    xnor g21003 ( n19360 , n2672 , n24567 );
    not g21004 ( n12450 , n11992 );
    xnor g21005 ( n18446 , n4093 , n2956 );
    not g21006 ( n9829 , n2024 );
    and g21007 ( n24534 , n6538 , n28362 );
    and g21008 ( n5526 , n2757 , n17995 );
    not g21009 ( n27682 , n7427 );
    not g21010 ( n16274 , n6858 );
    nor g21011 ( n20612 , n15363 , n4946 );
    nor g21012 ( n20615 , n2360 , n27532 );
    not g21013 ( n28658 , n11694 );
    not g21014 ( n19006 , n29667 );
    nor g21015 ( n3452 , n15413 , n14162 );
    or g21016 ( n28468 , n20030 , n7319 );
    or g21017 ( n12578 , n19221 , n6822 );
    and g21018 ( n1658 , n17045 , n17384 );
    and g21019 ( n11191 , n7245 , n22957 );
    and g21020 ( n20256 , n28551 , n28694 );
    or g21021 ( n7332 , n30840 , n5925 );
    xnor g21022 ( n28612 , n19066 , n19516 );
    nor g21023 ( n31714 , n16383 , n14080 );
    and g21024 ( n18935 , n711 , n30528 );
    nor g21025 ( n19500 , n31917 , n28489 );
    not g21026 ( n20111 , n20888 );
    or g21027 ( n10491 , n16008 , n28569 );
    xnor g21028 ( n1525 , n17428 , n24129 );
    xnor g21029 ( n12378 , n11443 , n24610 );
    not g21030 ( n6703 , n2603 );
    not g21031 ( n17563 , n9370 );
    xnor g21032 ( n1883 , n31455 , n10451 );
    not g21033 ( n11424 , n7770 );
    not g21034 ( n18783 , n18135 );
    or g21035 ( n18906 , n4927 , n25342 );
    not g21036 ( n11002 , n22367 );
    xnor g21037 ( n22114 , n29687 , n12317 );
    not g21038 ( n19583 , n27367 );
    or g21039 ( n31777 , n4469 , n18897 );
    not g21040 ( n12084 , n9026 );
    or g21041 ( n9442 , n16657 , n11207 );
    or g21042 ( n26039 , n2607 , n12738 );
    not g21043 ( n17813 , n13859 );
    or g21044 ( n14739 , n19559 , n20117 );
    and g21045 ( n13082 , n18023 , n15579 );
    or g21046 ( n22191 , n7780 , n16363 );
    xnor g21047 ( n18861 , n20299 , n4882 );
    xnor g21048 ( n21605 , n12642 , n30085 );
    and g21049 ( n27766 , n8303 , n26513 );
    xnor g21050 ( n14565 , n20903 , n13424 );
    and g21051 ( n12755 , n29730 , n29610 );
    or g21052 ( n21040 , n21026 , n17276 );
    or g21053 ( n17476 , n14520 , n12043 );
    nor g21054 ( n27299 , n2939 , n2231 );
    not g21055 ( n1685 , n17072 );
    not g21056 ( n184 , n22512 );
    or g21057 ( n3456 , n15069 , n17349 );
    and g21058 ( n25973 , n5507 , n22782 );
    or g21059 ( n29925 , n25084 , n19909 );
    not g21060 ( n8807 , n621 );
    and g21061 ( n10267 , n30108 , n2486 );
    or g21062 ( n10428 , n8024 , n5841 );
    or g21063 ( n31532 , n11802 , n30712 );
    or g21064 ( n26789 , n12676 , n5977 );
    xnor g21065 ( n2253 , n28925 , n18372 );
    xnor g21066 ( n3062 , n8635 , n30929 );
    or g21067 ( n5519 , n20236 , n11166 );
    or g21068 ( n6886 , n19374 , n6958 );
    xnor g21069 ( n25490 , n8834 , n10981 );
    xnor g21070 ( n27069 , n1996 , n18682 );
    xnor g21071 ( n6517 , n9877 , n11313 );
    xnor g21072 ( n1629 , n10492 , n788 );
    or g21073 ( n9833 , n24137 , n10302 );
    not g21074 ( n7274 , n20686 );
    not g21075 ( n4221 , n26387 );
    and g21076 ( n20033 , n8709 , n27371 );
    and g21077 ( n31130 , n28469 , n5235 );
    xnor g21078 ( n30710 , n11998 , n26636 );
    xnor g21079 ( n17957 , n7642 , n24464 );
    or g21080 ( n28333 , n2716 , n30322 );
    not g21081 ( n24097 , n9924 );
    or g21082 ( n23526 , n14908 , n21061 );
    or g21083 ( n9534 , n13335 , n25835 );
    not g21084 ( n8480 , n9177 );
    or g21085 ( n31430 , n11408 , n10743 );
    and g21086 ( n24566 , n13199 , n22231 );
    or g21087 ( n1625 , n22045 , n5132 );
    not g21088 ( n15036 , n11203 );
    buf g21089 ( n13554 , n10148 );
    or g21090 ( n22322 , n15833 , n31595 );
    nor g21091 ( n3264 , n9617 , n13272 );
    or g21092 ( n17453 , n27677 , n3137 );
    xnor g21093 ( n13158 , n23405 , n22504 );
    or g21094 ( n7448 , n10409 , n14607 );
    and g21095 ( n408 , n29222 , n25784 );
    xnor g21096 ( n28746 , n7224 , n22248 );
    nor g21097 ( n26028 , n25527 , n27453 );
    or g21098 ( n12843 , n12015 , n23059 );
    xnor g21099 ( n7992 , n16154 , n21673 );
    not g21100 ( n9600 , n23498 );
    not g21101 ( n10939 , n24890 );
    not g21102 ( n21327 , n29741 );
    not g21103 ( n109 , n13973 );
    xnor g21104 ( n12718 , n11710 , n31470 );
    not g21105 ( n19920 , n25626 );
    xnor g21106 ( n8213 , n4844 , n19538 );
    xnor g21107 ( n20718 , n5327 , n11168 );
    and g21108 ( n23865 , n18697 , n20325 );
    not g21109 ( n18082 , n25496 );
    xnor g21110 ( n17946 , n11040 , n7394 );
    not g21111 ( n13632 , n7986 );
    xnor g21112 ( n17943 , n18016 , n1420 );
    xnor g21113 ( n3516 , n12432 , n24558 );
    xnor g21114 ( n26319 , n13041 , n9358 );
    xnor g21115 ( n4621 , n23999 , n3593 );
    and g21116 ( n21948 , n1333 , n5792 );
    and g21117 ( n22400 , n31576 , n19781 );
    not g21118 ( n28600 , n23522 );
    or g21119 ( n2996 , n5770 , n10928 );
    or g21120 ( n15705 , n26369 , n8911 );
    xor g21121 ( n4361 , n5577 , n5897 );
    and g21122 ( n13371 , n16738 , n15637 );
    not g21123 ( n31914 , n7191 );
    and g21124 ( n24450 , n15575 , n3356 );
    and g21125 ( n20204 , n1826 , n30325 );
    or g21126 ( n19713 , n8521 , n435 );
    not g21127 ( n6068 , n8873 );
    and g21128 ( n3988 , n11669 , n6287 );
    or g21129 ( n28122 , n7760 , n10689 );
    not g21130 ( n16767 , n18830 );
    not g21131 ( n27292 , n18203 );
    xnor g21132 ( n22864 , n27802 , n23262 );
    or g21133 ( n17482 , n3582 , n27092 );
    xnor g21134 ( n20616 , n2942 , n23320 );
    or g21135 ( n12528 , n10818 , n14892 );
    not g21136 ( n10751 , n4844 );
    xnor g21137 ( n18639 , n6534 , n3108 );
    nor g21138 ( n309 , n3725 , n30843 );
    and g21139 ( n13924 , n619 , n24740 );
    not g21140 ( n20902 , n31426 );
    xnor g21141 ( n29885 , n2000 , n13975 );
    not g21142 ( n10123 , n16741 );
    nor g21143 ( n29284 , n24289 , n21661 );
    or g21144 ( n16323 , n1026 , n19893 );
    not g21145 ( n3926 , n17824 );
    xnor g21146 ( n5418 , n21972 , n23435 );
    not g21147 ( n26469 , n4523 );
    or g21148 ( n9819 , n18011 , n4137 );
    nor g21149 ( n21795 , n18759 , n10762 );
    xnor g21150 ( n9122 , n3152 , n11782 );
    not g21151 ( n31543 , n18114 );
    and g21152 ( n29124 , n14803 , n3109 );
    or g21153 ( n659 , n10112 , n14465 );
    or g21154 ( n20206 , n870 , n23466 );
    and g21155 ( n4066 , n21845 , n5513 );
    not g21156 ( n26168 , n16149 );
    or g21157 ( n28028 , n3174 , n22559 );
    not g21158 ( n10464 , n8948 );
    nor g21159 ( n31562 , n11626 , n1018 );
    not g21160 ( n22366 , n25369 );
    not g21161 ( n29632 , n31970 );
    or g21162 ( n1569 , n23494 , n26905 );
    or g21163 ( n20919 , n3259 , n13172 );
    or g21164 ( n3435 , n15922 , n1134 );
    and g21165 ( n7281 , n7572 , n19819 );
    not g21166 ( n23349 , n28267 );
    xor g21167 ( n29595 , n29855 , n31366 );
    xnor g21168 ( n25538 , n8931 , n15342 );
    and g21169 ( n15625 , n6811 , n9336 );
    xnor g21170 ( n11217 , n22870 , n8097 );
    or g21171 ( n29327 , n19550 , n30547 );
    or g21172 ( n13900 , n8447 , n1190 );
    xnor g21173 ( n14466 , n10747 , n11132 );
    xnor g21174 ( n13693 , n9201 , n18131 );
    xnor g21175 ( n20235 , n13604 , n1635 );
    nor g21176 ( n18490 , n30087 , n1328 );
    nor g21177 ( n8068 , n22145 , n12717 );
    not g21178 ( n25027 , n18660 );
    nor g21179 ( n15307 , n15436 , n10131 );
    xnor g21180 ( n7706 , n16810 , n13701 );
    xnor g21181 ( n15261 , n28157 , n26752 );
    nor g21182 ( n26898 , n24382 , n29520 );
    xnor g21183 ( n14580 , n26148 , n775 );
    or g21184 ( n22491 , n3001 , n12656 );
    and g21185 ( n22711 , n20209 , n107 );
    or g21186 ( n23200 , n13298 , n17244 );
    and g21187 ( n11490 , n24097 , n17910 );
    not g21188 ( n31688 , n20897 );
    not g21189 ( n1152 , n18221 );
    and g21190 ( n7555 , n4042 , n23322 );
    and g21191 ( n22561 , n6047 , n21880 );
    not g21192 ( n7459 , n28858 );
    not g21193 ( n15828 , n16882 );
    xnor g21194 ( n23970 , n18491 , n19733 );
    or g21195 ( n17892 , n21871 , n1915 );
    xnor g21196 ( n29762 , n15401 , n23643 );
    or g21197 ( n9937 , n19405 , n17339 );
    or g21198 ( n11742 , n10311 , n14943 );
    or g21199 ( n24172 , n13334 , n8646 );
    xnor g21200 ( n17040 , n1652 , n14363 );
    not g21201 ( n3299 , n3261 );
    and g21202 ( n14532 , n5547 , n9292 );
    and g21203 ( n21546 , n12621 , n1616 );
    or g21204 ( n17804 , n24893 , n25374 );
    and g21205 ( n29185 , n17216 , n8133 );
    xnor g21206 ( n26483 , n15579 , n18023 );
    or g21207 ( n25286 , n724 , n17124 );
    nor g21208 ( n4142 , n2592 , n26481 );
    not g21209 ( n20056 , n10264 );
    or g21210 ( n1599 , n12629 , n15623 );
    xnor g21211 ( n6260 , n27036 , n15265 );
    xnor g21212 ( n2165 , n22879 , n5893 );
    or g21213 ( n24752 , n21493 , n20917 );
    xnor g21214 ( n12678 , n7195 , n22138 );
    xnor g21215 ( n16426 , n16674 , n11462 );
    or g21216 ( n2751 , n15377 , n748 );
    or g21217 ( n9916 , n14617 , n31695 );
    not g21218 ( n3883 , n12777 );
    xnor g21219 ( n8699 , n30245 , n12566 );
    xnor g21220 ( n22719 , n27077 , n12207 );
    nor g21221 ( n13008 , n29642 , n29836 );
    and g21222 ( n6379 , n25302 , n10771 );
    xnor g21223 ( n26400 , n22423 , n12035 );
    not g21224 ( n25669 , n26181 );
    xnor g21225 ( n5965 , n5277 , n6372 );
    not g21226 ( n1490 , n28268 );
    or g21227 ( n13561 , n15633 , n415 );
    nor g21228 ( n25605 , n30908 , n21055 );
    xnor g21229 ( n25487 , n6288 , n17386 );
    xnor g21230 ( n28306 , n4692 , n1554 );
    or g21231 ( n24367 , n22487 , n27402 );
    not g21232 ( n251 , n26507 );
    not g21233 ( n4425 , n28006 );
    and g21234 ( n9103 , n24637 , n29093 );
    not g21235 ( n60 , n2968 );
    and g21236 ( n30576 , n8609 , n1337 );
    xnor g21237 ( n8253 , n1340 , n5144 );
    nor g21238 ( n294 , n19132 , n15604 );
    not g21239 ( n387 , n27148 );
    xnor g21240 ( n20808 , n22448 , n21783 );
    or g21241 ( n1470 , n25478 , n5198 );
    not g21242 ( n28937 , n14942 );
    or g21243 ( n25965 , n20865 , n12183 );
    not g21244 ( n11523 , n11121 );
    not g21245 ( n25670 , n6338 );
    not g21246 ( n24574 , n20270 );
    or g21247 ( n3300 , n23251 , n2376 );
    xnor g21248 ( n23416 , n26468 , n7308 );
    and g21249 ( n20738 , n2445 , n505 );
    or g21250 ( n28373 , n15896 , n14299 );
    or g21251 ( n19284 , n10562 , n25013 );
    not g21252 ( n1293 , n929 );
    nor g21253 ( n27580 , n30203 , n15039 );
    nor g21254 ( n20970 , n15427 , n19445 );
    xnor g21255 ( n3791 , n9523 , n4757 );
    nor g21256 ( n30861 , n17948 , n29336 );
    xnor g21257 ( n1550 , n9701 , n14231 );
    nor g21258 ( n19962 , n9336 , n1675 );
    not g21259 ( n23410 , n18527 );
    xnor g21260 ( n7265 , n25634 , n7899 );
    nor g21261 ( n26983 , n26339 , n17040 );
    not g21262 ( n8934 , n2244 );
    not g21263 ( n5775 , n7413 );
    or g21264 ( n17676 , n20700 , n8618 );
    xnor g21265 ( n12454 , n12236 , n30489 );
    and g21266 ( n5787 , n3866 , n24867 );
    xor g21267 ( n5025 , n22139 , n19615 );
    xnor g21268 ( n31408 , n30314 , n2975 );
    not g21269 ( n19563 , n13079 );
    or g21270 ( n15330 , n8972 , n15460 );
    not g21271 ( n11414 , n12031 );
    or g21272 ( n13362 , n24455 , n29721 );
    nor g21273 ( n7584 , n3471 , n6040 );
    and g21274 ( n17844 , n30995 , n5486 );
    not g21275 ( n26485 , n29120 );
    and g21276 ( n9911 , n31154 , n3751 );
    or g21277 ( n4442 , n31019 , n73 );
    and g21278 ( n12056 , n12235 , n15881 );
    not g21279 ( n25765 , n29436 );
    not g21280 ( n7489 , n17533 );
    nor g21281 ( n18061 , n20625 , n31754 );
    nor g21282 ( n17366 , n12762 , n12619 );
    or g21283 ( n3903 , n25368 , n5520 );
    and g21284 ( n15343 , n5542 , n21363 );
    nor g21285 ( n8425 , n6349 , n22279 );
    not g21286 ( n1777 , n11387 );
    or g21287 ( n30628 , n16410 , n12351 );
    and g21288 ( n5887 , n5558 , n6196 );
    and g21289 ( n15189 , n706 , n19178 );
    or g21290 ( n27551 , n14742 , n4778 );
    xnor g21291 ( n15845 , n31674 , n28261 );
    not g21292 ( n23475 , n31085 );
    xnor g21293 ( n29918 , n30696 , n27830 );
    xnor g21294 ( n14205 , n26451 , n18918 );
    not g21295 ( n27704 , n24202 );
    xnor g21296 ( n30338 , n21983 , n6700 );
    not g21297 ( n1955 , n6507 );
    xnor g21298 ( n3172 , n8993 , n31115 );
    nor g21299 ( n9736 , n20453 , n30769 );
    xnor g21300 ( n8402 , n29249 , n2231 );
    xnor g21301 ( n16623 , n24188 , n23555 );
    or g21302 ( n25293 , n3859 , n30663 );
    xnor g21303 ( n7938 , n27738 , n20891 );
    and g21304 ( n7132 , n15344 , n4989 );
    and g21305 ( n26938 , n12885 , n19634 );
    not g21306 ( n17046 , n7967 );
    xnor g21307 ( n7485 , n30070 , n10994 );
    xnor g21308 ( n28691 , n7892 , n6626 );
    xnor g21309 ( n17495 , n6120 , n21772 );
    or g21310 ( n26360 , n8062 , n18956 );
    xnor g21311 ( n13688 , n5821 , n20320 );
    xnor g21312 ( n32018 , n26648 , n3415 );
    and g21313 ( n10617 , n22771 , n28016 );
    xnor g21314 ( n31215 , n2041 , n30411 );
    not g21315 ( n14861 , n28230 );
    not g21316 ( n4070 , n6502 );
    nor g21317 ( n11018 , n12411 , n13352 );
    or g21318 ( n19242 , n5314 , n17213 );
    and g21319 ( n83 , n31300 , n30288 );
    and g21320 ( n16874 , n18273 , n30011 );
    not g21321 ( n6569 , n14227 );
    or g21322 ( n16611 , n22886 , n12856 );
    and g21323 ( n30879 , n10481 , n11091 );
    xnor g21324 ( n14716 , n31154 , n29266 );
    or g21325 ( n21991 , n5502 , n10642 );
    or g21326 ( n9247 , n23422 , n5997 );
    xnor g21327 ( n19051 , n25352 , n30503 );
    xor g21328 ( n25546 , n8830 , n24251 );
    and g21329 ( n5970 , n16265 , n8230 );
    xnor g21330 ( n23489 , n1819 , n13494 );
    not g21331 ( n24527 , n11080 );
    or g21332 ( n28137 , n19522 , n10285 );
    or g21333 ( n2472 , n10716 , n2054 );
    and g21334 ( n18885 , n21022 , n16949 );
    xnor g21335 ( n10879 , n20333 , n30709 );
    or g21336 ( n29299 , n11490 , n26209 );
    xnor g21337 ( n3439 , n12543 , n15245 );
    xor g21338 ( n28170 , n26102 , n5313 );
    xnor g21339 ( n28872 , n5005 , n13479 );
    and g21340 ( n16684 , n8040 , n23209 );
    xnor g21341 ( n20260 , n31839 , n5838 );
    or g21342 ( n21005 , n4500 , n27746 );
    buf g21343 ( n27089 , n20998 );
    or g21344 ( n15601 , n3993 , n5209 );
    nor g21345 ( n26380 , n16560 , n16259 );
    not g21346 ( n17115 , n7128 );
    or g21347 ( n19253 , n19532 , n25459 );
    or g21348 ( n19866 , n6527 , n27379 );
    xnor g21349 ( n31878 , n24027 , n25178 );
    or g21350 ( n5872 , n19840 , n15333 );
    nor g21351 ( n26841 , n7718 , n16934 );
    and g21352 ( n16343 , n27529 , n23269 );
    not g21353 ( n5358 , n6789 );
    not g21354 ( n12283 , n22577 );
    not g21355 ( n19408 , n18623 );
    nor g21356 ( n31006 , n22922 , n20474 );
    or g21357 ( n23457 , n9269 , n1425 );
    xnor g21358 ( n9540 , n31668 , n26961 );
    not g21359 ( n2627 , n29840 );
    and g21360 ( n7573 , n5564 , n5181 );
    or g21361 ( n19833 , n1879 , n21393 );
    nor g21362 ( n11909 , n4541 , n9611 );
    xnor g21363 ( n14378 , n25340 , n15476 );
    nor g21364 ( n2087 , n14598 , n27368 );
    xnor g21365 ( n29980 , n31203 , n22587 );
    not g21366 ( n16456 , n18497 );
    not g21367 ( n27859 , n18919 );
    xnor g21368 ( n11272 , n11533 , n30669 );
    and g21369 ( n17714 , n31274 , n1993 );
    xnor g21370 ( n1785 , n10160 , n5446 );
    xnor g21371 ( n15334 , n25402 , n2798 );
    not g21372 ( n6232 , n19217 );
    and g21373 ( n4010 , n12483 , n12239 );
    or g21374 ( n15033 , n30570 , n20638 );
    not g21375 ( n11478 , n20390 );
    or g21376 ( n16176 , n9726 , n6928 );
    not g21377 ( n13845 , n16369 );
    xnor g21378 ( n9733 , n27217 , n18381 );
    and g21379 ( n20008 , n25668 , n6803 );
    not g21380 ( n5763 , n22396 );
    and g21381 ( n10462 , n4792 , n219 );
    xnor g21382 ( n1761 , n8156 , n23869 );
    and g21383 ( n15739 , n23660 , n8407 );
    xnor g21384 ( n4158 , n22239 , n22931 );
    xnor g21385 ( n9010 , n26423 , n12979 );
    not g21386 ( n3363 , n14641 );
    not g21387 ( n12266 , n27975 );
    xnor g21388 ( n29041 , n28081 , n15999 );
    nor g21389 ( n27180 , n25954 , n2748 );
    or g21390 ( n2863 , n31918 , n8579 );
    not g21391 ( n5428 , n8824 );
    or g21392 ( n14971 , n2912 , n239 );
    not g21393 ( n31764 , n27384 );
    or g21394 ( n3601 , n30610 , n13095 );
    or g21395 ( n7405 , n5831 , n19720 );
    xnor g21396 ( n26599 , n3837 , n24086 );
    xnor g21397 ( n19670 , n14498 , n18669 );
    not g21398 ( n18272 , n21024 );
    not g21399 ( n10669 , n17762 );
    and g21400 ( n11741 , n1922 , n6793 );
    or g21401 ( n6410 , n3266 , n10815 );
    xnor g21402 ( n9317 , n31256 , n7605 );
    xnor g21403 ( n9077 , n27012 , n3326 );
    not g21404 ( n25434 , n17447 );
    not g21405 ( n31516 , n27783 );
    nor g21406 ( n22099 , n10598 , n31078 );
    not g21407 ( n12955 , n16314 );
    xnor g21408 ( n14323 , n3599 , n11253 );
    and g21409 ( n4449 , n28359 , n21156 );
    buf g21410 ( n26496 , n23968 );
    not g21411 ( n5384 , n8252 );
    nor g21412 ( n16242 , n11677 , n31603 );
    not g21413 ( n15408 , n20627 );
    or g21414 ( n4392 , n15699 , n22291 );
    not g21415 ( n13038 , n20786 );
    not g21416 ( n13716 , n1307 );
    xor g21417 ( n17901 , n11440 , n3907 );
    and g21418 ( n15597 , n25815 , n25100 );
    or g21419 ( n168 , n8361 , n10634 );
    xnor g21420 ( n14786 , n26172 , n276 );
    or g21421 ( n27363 , n10227 , n14253 );
    not g21422 ( n16088 , n28786 );
    not g21423 ( n15897 , n24918 );
    and g21424 ( n7499 , n12021 , n22535 );
    or g21425 ( n7846 , n8464 , n7555 );
    xnor g21426 ( n20589 , n8148 , n18508 );
    xnor g21427 ( n3630 , n10152 , n24568 );
    xnor g21428 ( n14685 , n10428 , n5080 );
    not g21429 ( n10598 , n30201 );
    xnor g21430 ( n24570 , n10027 , n13266 );
    nor g21431 ( n24978 , n22316 , n21466 );
    nor g21432 ( n19401 , n27896 , n10734 );
    not g21433 ( n18920 , n1680 );
    and g21434 ( n28777 , n15676 , n4662 );
    or g21435 ( n4655 , n8376 , n25243 );
    xnor g21436 ( n10163 , n9537 , n19066 );
    or g21437 ( n27324 , n1756 , n19813 );
    not g21438 ( n15433 , n19177 );
    nor g21439 ( n24234 , n24970 , n11313 );
    and g21440 ( n19585 , n23243 , n8002 );
    or g21441 ( n14881 , n27208 , n4036 );
    not g21442 ( n22994 , n21111 );
    not g21443 ( n12299 , n25682 );
    not g21444 ( n14943 , n3802 );
    not g21445 ( n28061 , n30232 );
    and g21446 ( n4908 , n15651 , n13779 );
    and g21447 ( n10970 , n19191 , n7536 );
    not g21448 ( n23171 , n15522 );
    not g21449 ( n18979 , n20101 );
    xnor g21450 ( n21421 , n7079 , n13912 );
    and g21451 ( n5540 , n1440 , n25441 );
    xnor g21452 ( n20716 , n20344 , n19406 );
    not g21453 ( n21020 , n23840 );
    not g21454 ( n29441 , n10989 );
    nor g21455 ( n17201 , n5964 , n6247 );
    xnor g21456 ( n3274 , n3111 , n31866 );
    or g21457 ( n21088 , n8008 , n30258 );
    and g21458 ( n21027 , n1463 , n1482 );
    or g21459 ( n17307 , n4850 , n9698 );
    or g21460 ( n7509 , n24008 , n5716 );
    xnor g21461 ( n30723 , n282 , n26956 );
    not g21462 ( n5612 , n11815 );
    xnor g21463 ( n12495 , n3137 , n28746 );
    nor g21464 ( n6067 , n4424 , n4757 );
    and g21465 ( n8299 , n24239 , n17118 );
    xnor g21466 ( n2113 , n28468 , n592 );
    xnor g21467 ( n27689 , n18398 , n30852 );
    or g21468 ( n16738 , n12891 , n23132 );
    or g21469 ( n26230 , n24297 , n16996 );
    xnor g21470 ( n28095 , n8877 , n20549 );
    not g21471 ( n7642 , n2410 );
    xnor g21472 ( n15570 , n1426 , n15215 );
    xnor g21473 ( n28491 , n13397 , n23648 );
    or g21474 ( n10386 , n17211 , n8697 );
    not g21475 ( n11121 , n13934 );
    xnor g21476 ( n11996 , n16299 , n891 );
    and g21477 ( n16829 , n6903 , n18909 );
    xnor g21478 ( n31709 , n18615 , n27226 );
    nor g21479 ( n18547 , n29141 , n27758 );
    xnor g21480 ( n21006 , n25291 , n7184 );
    and g21481 ( n2406 , n22448 , n19277 );
    nor g21482 ( n29563 , n22706 , n31253 );
    not g21483 ( n5616 , n404 );
    xnor g21484 ( n13065 , n21522 , n15749 );
    and g21485 ( n26557 , n6145 , n26923 );
    not g21486 ( n13089 , n13011 );
    and g21487 ( n1661 , n18970 , n21005 );
    xor g21488 ( n10630 , n21871 , n19810 );
    not g21489 ( n27487 , n7396 );
    not g21490 ( n23867 , n27884 );
    not g21491 ( n22053 , n416 );
    or g21492 ( n28082 , n5627 , n9981 );
    not g21493 ( n30862 , n18832 );
    xnor g21494 ( n4225 , n10158 , n23561 );
    not g21495 ( n27791 , n1710 );
    xnor g21496 ( n1783 , n4189 , n2275 );
    or g21497 ( n8501 , n18411 , n26048 );
    not g21498 ( n3335 , n5683 );
    not g21499 ( n18930 , n7004 );
    xnor g21500 ( n6021 , n26324 , n31050 );
    xnor g21501 ( n1562 , n7353 , n3244 );
    or g21502 ( n18031 , n17496 , n22416 );
    not g21503 ( n5188 , n4488 );
    not g21504 ( n26931 , n10357 );
    nor g21505 ( n619 , n5355 , n7874 );
    not g21506 ( n19000 , n17653 );
    and g21507 ( n15180 , n19047 , n16226 );
    or g21508 ( n28994 , n25188 , n7710 );
    or g21509 ( n20610 , n27192 , n12693 );
    xnor g21510 ( n26056 , n24132 , n2483 );
    xnor g21511 ( n10156 , n22537 , n26980 );
    and g21512 ( n27415 , n4945 , n25799 );
    not g21513 ( n13935 , n11253 );
    not g21514 ( n25570 , n10443 );
    xnor g21515 ( n4287 , n1454 , n21185 );
    or g21516 ( n19341 , n25403 , n26555 );
    xnor g21517 ( n31650 , n2852 , n28225 );
    and g21518 ( n28567 , n30638 , n11532 );
    or g21519 ( n12088 , n5388 , n16847 );
    xnor g21520 ( n8456 , n27488 , n21307 );
    and g21521 ( n28196 , n1390 , n5644 );
    xnor g21522 ( n22832 , n16065 , n24781 );
    xor g21523 ( n27865 , n8065 , n1924 );
    and g21524 ( n20849 , n29485 , n3164 );
    xnor g21525 ( n17470 , n10616 , n10511 );
    not g21526 ( n28087 , n23043 );
    or g21527 ( n28631 , n5767 , n20378 );
    nor g21528 ( n10628 , n25827 , n23991 );
    xor g21529 ( n20109 , n15854 , n671 );
    or g21530 ( n9226 , n15407 , n1731 );
    xnor g21531 ( n28989 , n22725 , n11725 );
    xnor g21532 ( n6307 , n16747 , n2231 );
    or g21533 ( n25909 , n30273 , n29710 );
    or g21534 ( n10360 , n12712 , n7055 );
    buf g21535 ( n31146 , n20813 );
    or g21536 ( n24108 , n8425 , n6214 );
    or g21537 ( n18965 , n18067 , n22104 );
    and g21538 ( n26475 , n27296 , n29511 );
    and g21539 ( n6065 , n13339 , n23 );
    not g21540 ( n2920 , n11962 );
    xnor g21541 ( n11023 , n12866 , n20703 );
    not g21542 ( n19393 , n21743 );
    or g21543 ( n24559 , n28981 , n19077 );
    or g21544 ( n3823 , n14850 , n24497 );
    or g21545 ( n20741 , n974 , n23775 );
    not g21546 ( n12918 , n30271 );
    and g21547 ( n28059 , n18215 , n12714 );
    and g21548 ( n2198 , n20688 , n18043 );
    nor g21549 ( n14168 , n24128 , n395 );
    xnor g21550 ( n31171 , n11262 , n22434 );
    and g21551 ( n19547 , n67 , n31746 );
    nor g21552 ( n23990 , n30179 , n15169 );
    or g21553 ( n7250 , n17740 , n10265 );
    xnor g21554 ( n14546 , n30154 , n17053 );
    or g21555 ( n20884 , n14496 , n11916 );
    xnor g21556 ( n29736 , n21574 , n11242 );
    not g21557 ( n25078 , n20837 );
    and g21558 ( n1454 , n25402 , n23932 );
    xnor g21559 ( n18469 , n31320 , n31539 );
    and g21560 ( n10246 , n6847 , n13722 );
    not g21561 ( n18841 , n24712 );
    not g21562 ( n11826 , n24834 );
    or g21563 ( n15911 , n31918 , n28306 );
    or g21564 ( n19996 , n5538 , n21797 );
    and g21565 ( n4948 , n19072 , n7383 );
    xnor g21566 ( n13374 , n22046 , n12467 );
    xnor g21567 ( n6489 , n11173 , n1784 );
    nor g21568 ( n18028 , n28574 , n13492 );
    and g21569 ( n10780 , n13464 , n23554 );
    xnor g21570 ( n7179 , n29728 , n1815 );
    nor g21571 ( n10062 , n3036 , n4812 );
    not g21572 ( n13543 , n12502 );
    or g21573 ( n5958 , n14813 , n21565 );
    or g21574 ( n17725 , n30515 , n25029 );
    not g21575 ( n21034 , n2997 );
    not g21576 ( n29056 , n31853 );
    xnor g21577 ( n1265 , n23713 , n13118 );
    or g21578 ( n15893 , n17026 , n12979 );
    xnor g21579 ( n6442 , n15923 , n11471 );
    and g21580 ( n12585 , n4615 , n26408 );
    or g21581 ( n1339 , n20905 , n23959 );
    and g21582 ( n26873 , n30033 , n7919 );
    xnor g21583 ( n26425 , n24855 , n3585 );
    or g21584 ( n3517 , n6434 , n15562 );
    or g21585 ( n26127 , n23563 , n28585 );
    xnor g21586 ( n23398 , n17576 , n10723 );
    not g21587 ( n7408 , n15191 );
    xnor g21588 ( n15107 , n16587 , n31182 );
    nor g21589 ( n18576 , n24081 , n12048 );
    or g21590 ( n2474 , n17014 , n6522 );
    or g21591 ( n29275 , n19825 , n26810 );
    not g21592 ( n4776 , n20510 );
    or g21593 ( n17961 , n30044 , n12202 );
    and g21594 ( n12836 , n24801 , n16907 );
    or g21595 ( n25839 , n31168 , n9859 );
    not g21596 ( n12880 , n19224 );
    xnor g21597 ( n4967 , n4253 , n31889 );
    not g21598 ( n28293 , n9691 );
    or g21599 ( n2314 , n405 , n25766 );
    or g21600 ( n25725 , n15992 , n25594 );
    nor g21601 ( n18132 , n18667 , n26082 );
    xnor g21602 ( n959 , n30550 , n28832 );
    or g21603 ( n18383 , n10142 , n1672 );
    not g21604 ( n20924 , n23701 );
    or g21605 ( n6996 , n16609 , n29568 );
    nor g21606 ( n16311 , n13140 , n19155 );
    nor g21607 ( n7242 , n2298 , n5081 );
    not g21608 ( n7566 , n17227 );
    and g21609 ( n21016 , n14048 , n8719 );
    or g21610 ( n11383 , n1163 , n24592 );
    or g21611 ( n26986 , n7216 , n13318 );
    not g21612 ( n12540 , n19033 );
    and g21613 ( n4712 , n25140 , n23679 );
    xnor g21614 ( n28507 , n15461 , n5942 );
    or g21615 ( n6289 , n11486 , n1435 );
    nor g21616 ( n2713 , n25793 , n7127 );
    xnor g21617 ( n1892 , n664 , n14690 );
    xnor g21618 ( n3002 , n12581 , n1501 );
    or g21619 ( n9707 , n10566 , n13909 );
    or g21620 ( n14840 , n149 , n23234 );
    or g21621 ( n30127 , n16295 , n10573 );
    not g21622 ( n1442 , n7193 );
    xnor g21623 ( n25620 , n24462 , n2059 );
    not g21624 ( n31698 , n20020 );
    and g21625 ( n19825 , n2430 , n26207 );
    or g21626 ( n5127 , n28411 , n26337 );
    nor g21627 ( n5530 , n8931 , n26889 );
    or g21628 ( n22918 , n21289 , n3564 );
    not g21629 ( n25206 , n1048 );
    xnor g21630 ( n5517 , n11230 , n17604 );
    or g21631 ( n11817 , n13607 , n5700 );
    xnor g21632 ( n15364 , n22644 , n19517 );
    and g21633 ( n16542 , n10613 , n12876 );
    not g21634 ( n29288 , n20343 );
    not g21635 ( n27266 , n18657 );
    or g21636 ( n23346 , n13366 , n17555 );
    or g21637 ( n31291 , n11645 , n13948 );
    xnor g21638 ( n8600 , n2879 , n3281 );
    and g21639 ( n9735 , n12915 , n28163 );
    xnor g21640 ( n16608 , n3742 , n17875 );
    not g21641 ( n10085 , n21466 );
    and g21642 ( n12387 , n15072 , n30430 );
    xnor g21643 ( n2375 , n30617 , n7131 );
    and g21644 ( n17848 , n21501 , n13581 );
    and g21645 ( n22876 , n27395 , n25671 );
    and g21646 ( n3098 , n5311 , n30350 );
    not g21647 ( n9850 , n31448 );
    not g21648 ( n818 , n13148 );
    or g21649 ( n24553 , n3907 , n11345 );
    not g21650 ( n20898 , n29824 );
    nor g21651 ( n20521 , n1139 , n13083 );
    not g21652 ( n13516 , n30843 );
    not g21653 ( n3364 , n20554 );
    and g21654 ( n14914 , n28090 , n19732 );
    nor g21655 ( n4207 , n11692 , n16525 );
    not g21656 ( n6393 , n15144 );
    xnor g21657 ( n31622 , n21489 , n8536 );
    xnor g21658 ( n5226 , n16353 , n27553 );
    and g21659 ( n8116 , n26304 , n27987 );
    not g21660 ( n22058 , n29439 );
    or g21661 ( n1611 , n27995 , n14368 );
    or g21662 ( n20778 , n15376 , n2289 );
    not g21663 ( n10218 , n8764 );
    and g21664 ( n9713 , n23747 , n12395 );
    or g21665 ( n7991 , n3108 , n30822 );
    or g21666 ( n24374 , n18000 , n352 );
    not g21667 ( n30203 , n28209 );
    not g21668 ( n31438 , n5485 );
    not g21669 ( n4928 , n5047 );
    and g21670 ( n19009 , n24428 , n2390 );
    and g21671 ( n10530 , n13970 , n9189 );
    or g21672 ( n21691 , n13274 , n23315 );
    not g21673 ( n4822 , n12674 );
    not g21674 ( n6327 , n17536 );
    or g21675 ( n27283 , n1199 , n12486 );
    not g21676 ( n29787 , n15083 );
    xnor g21677 ( n23112 , n14244 , n27412 );
    xnor g21678 ( n18086 , n17724 , n7426 );
    not g21679 ( n6609 , n13640 );
    nor g21680 ( n1233 , n30425 , n17109 );
    nor g21681 ( n18338 , n31790 , n22746 );
    xnor g21682 ( n30257 , n20210 , n25758 );
    and g21683 ( n31133 , n26109 , n29801 );
    not g21684 ( n11964 , n19737 );
    xnor g21685 ( n17099 , n25334 , n4054 );
    nor g21686 ( n21567 , n31813 , n29121 );
    not g21687 ( n27200 , n9996 );
    xnor g21688 ( n30214 , n3076 , n20236 );
    and g21689 ( n17518 , n18076 , n19217 );
    xnor g21690 ( n29434 , n6822 , n19221 );
    or g21691 ( n27395 , n30576 , n10275 );
    not g21692 ( n18448 , n17833 );
    xnor g21693 ( n28325 , n6173 , n4720 );
    not g21694 ( n10151 , n28804 );
    not g21695 ( n12082 , n23187 );
    not g21696 ( n31100 , n4742 );
    not g21697 ( n24582 , n17844 );
    or g21698 ( n26057 , n1312 , n16352 );
    not g21699 ( n22319 , n18955 );
    buf g21700 ( n23597 , n8462 );
    not g21701 ( n12770 , n17793 );
    not g21702 ( n19125 , n2898 );
    nor g21703 ( n8637 , n21301 , n683 );
    not g21704 ( n17977 , n1980 );
    xnor g21705 ( n7478 , n19914 , n26302 );
    xnor g21706 ( n25037 , n31251 , n2608 );
    nor g21707 ( n13529 , n2438 , n31627 );
    or g21708 ( n7442 , n10060 , n1806 );
    and g21709 ( n1056 , n8441 , n22526 );
    xnor g21710 ( n8191 , n16990 , n11068 );
    not g21711 ( n9080 , n14492 );
    xnor g21712 ( n29761 , n940 , n5840 );
    xnor g21713 ( n10640 , n2867 , n25308 );
    and g21714 ( n18641 , n21775 , n11659 );
    or g21715 ( n22380 , n12881 , n5373 );
    not g21716 ( n5848 , n3025 );
    not g21717 ( n23348 , n2559 );
    or g21718 ( n19772 , n25145 , n23498 );
    xnor g21719 ( n22848 , n16821 , n27632 );
    or g21720 ( n16232 , n28629 , n16397 );
    not g21721 ( n28776 , n20050 );
    and g21722 ( n1151 , n931 , n614 );
    xnor g21723 ( n13767 , n27089 , n7209 );
    not g21724 ( n14025 , n7400 );
    xnor g21725 ( n10692 , n17276 , n31408 );
    not g21726 ( n31098 , n22981 );
    xnor g21727 ( n30713 , n27149 , n8915 );
    or g21728 ( n17071 , n4956 , n12295 );
    or g21729 ( n28534 , n154 , n11905 );
    buf g21730 ( n4571 , n10075 );
    nor g21731 ( n13631 , n23343 , n13387 );
    or g21732 ( n11914 , n18713 , n22435 );
    or g21733 ( n5196 , n3512 , n7625 );
    or g21734 ( n31712 , n28780 , n440 );
    not g21735 ( n14912 , n9275 );
    xnor g21736 ( n458 , n30386 , n5418 );
    or g21737 ( n7324 , n13381 , n31362 );
    buf g21738 ( n6717 , n22505 );
    and g21739 ( n25748 , n19281 , n20457 );
    and g21740 ( n1030 , n14936 , n12210 );
    or g21741 ( n9166 , n6414 , n12351 );
    xnor g21742 ( n24609 , n10071 , n25793 );
    not g21743 ( n15980 , n5290 );
    or g21744 ( n4805 , n15996 , n3115 );
    xnor g21745 ( n25543 , n21697 , n12799 );
    not g21746 ( n8316 , n14952 );
    or g21747 ( n11145 , n3432 , n31467 );
    not g21748 ( n2683 , n15010 );
    and g21749 ( n1795 , n29358 , n14810 );
    nor g21750 ( n13524 , n1125 , n10370 );
    not g21751 ( n27762 , n21581 );
    xor g21752 ( n16047 , n6293 , n17589 );
    or g21753 ( n5714 , n29737 , n4441 );
    not g21754 ( n22622 , n20774 );
    not g21755 ( n12851 , n24336 );
    and g21756 ( n3148 , n10754 , n31609 );
    or g21757 ( n7752 , n12580 , n988 );
    not g21758 ( n5567 , n21010 );
    xnor g21759 ( n20275 , n4926 , n26929 );
    nor g21760 ( n8371 , n12398 , n7028 );
    and g21761 ( n9294 , n21791 , n24359 );
    and g21762 ( n23690 , n27567 , n20415 );
    not g21763 ( n22997 , n4594 );
    and g21764 ( n29699 , n4893 , n6049 );
    not g21765 ( n4229 , n29591 );
    xnor g21766 ( n13681 , n2749 , n13137 );
    xnor g21767 ( n24943 , n12175 , n30201 );
    xnor g21768 ( n7710 , n10702 , n16471 );
    nor g21769 ( n19540 , n22233 , n5078 );
    or g21770 ( n12369 , n6870 , n29735 );
    not g21771 ( n11791 , n20627 );
    and g21772 ( n15480 , n16667 , n27797 );
    not g21773 ( n13509 , n22756 );
    not g21774 ( n9324 , n14624 );
    or g21775 ( n26472 , n20390 , n6787 );
    xnor g21776 ( n17387 , n26085 , n21050 );
    xnor g21777 ( n13657 , n9621 , n25700 );
    not g21778 ( n11321 , n11138 );
    xnor g21779 ( n18336 , n13469 , n20613 );
    or g21780 ( n22376 , n5387 , n2235 );
    xnor g21781 ( n20882 , n8309 , n25991 );
    not g21782 ( n6426 , n12072 );
    xnor g21783 ( n13933 , n14761 , n16441 );
    not g21784 ( n17882 , n4983 );
    and g21785 ( n27755 , n29882 , n18782 );
    or g21786 ( n13620 , n56 , n30484 );
    or g21787 ( n18187 , n1039 , n10474 );
    xnor g21788 ( n28205 , n16644 , n29630 );
    not g21789 ( n6191 , n31722 );
    or g21790 ( n29286 , n1111 , n29481 );
    nor g21791 ( n27653 , n10269 , n9455 );
    or g21792 ( n15982 , n4278 , n5543 );
    xnor g21793 ( n8672 , n31576 , n5231 );
    or g21794 ( n27576 , n12140 , n9339 );
    xnor g21795 ( n17041 , n19651 , n22123 );
    xnor g21796 ( n7285 , n27309 , n17844 );
    xnor g21797 ( n306 , n11789 , n6603 );
    xnor g21798 ( n11076 , n1178 , n9895 );
    and g21799 ( n27098 , n2822 , n11942 );
    not g21800 ( n19159 , n19312 );
    xnor g21801 ( n16980 , n3080 , n9591 );
    and g21802 ( n2401 , n8874 , n11051 );
    or g21803 ( n26937 , n3377 , n17430 );
    nor g21804 ( n18248 , n7009 , n18575 );
    xnor g21805 ( n232 , n554 , n256 );
    nor g21806 ( n8263 , n27453 , n24161 );
    or g21807 ( n7069 , n24814 , n30465 );
    or g21808 ( n27744 , n5069 , n11048 );
    not g21809 ( n17604 , n29559 );
    nor g21810 ( n26020 , n3307 , n20492 );
    not g21811 ( n26866 , n19632 );
    or g21812 ( n26499 , n23791 , n4762 );
    xnor g21813 ( n27839 , n1021 , n22390 );
    xnor g21814 ( n9860 , n15613 , n21310 );
    not g21815 ( n29574 , n25995 );
    xnor g21816 ( n15838 , n20166 , n26150 );
    not g21817 ( n25409 , n11193 );
    or g21818 ( n30748 , n27200 , n26931 );
    not g21819 ( n6340 , n11747 );
    or g21820 ( n11591 , n21105 , n24784 );
    and g21821 ( n29347 , n7892 , n6626 );
    xnor g21822 ( n29306 , n16698 , n30910 );
    or g21823 ( n1209 , n26177 , n8176 );
    not g21824 ( n27062 , n19752 );
    nor g21825 ( n8019 , n1346 , n17696 );
    not g21826 ( n14180 , n25872 );
    not g21827 ( n19339 , n15438 );
    xnor g21828 ( n15127 , n19128 , n13982 );
    or g21829 ( n28659 , n12172 , n20387 );
    xnor g21830 ( n9124 , n17881 , n24494 );
    or g21831 ( n9288 , n2546 , n23065 );
    xnor g21832 ( n16837 , n2887 , n808 );
    xnor g21833 ( n18379 , n4554 , n31889 );
    xnor g21834 ( n16096 , n12003 , n8239 );
    or g21835 ( n4136 , n28820 , n17846 );
    and g21836 ( n30460 , n10452 , n24867 );
    not g21837 ( n12145 , n11972 );
    nor g21838 ( n2835 , n16608 , n2864 );
    nor g21839 ( n16734 , n24601 , n9028 );
    not g21840 ( n37 , n4606 );
    not g21841 ( n19471 , n31519 );
    xnor g21842 ( n25757 , n30877 , n3522 );
    or g21843 ( n10827 , n16342 , n12825 );
    not g21844 ( n30418 , n6596 );
    not g21845 ( n18260 , n26961 );
    xnor g21846 ( n31733 , n11356 , n7921 );
    and g21847 ( n4581 , n26434 , n25081 );
    not g21848 ( n29571 , n25805 );
    xnor g21849 ( n31999 , n28010 , n23338 );
    nor g21850 ( n2098 , n12922 , n25695 );
    xnor g21851 ( n13256 , n17074 , n20067 );
    and g21852 ( n9737 , n7395 , n10388 );
    nor g21853 ( n1943 , n6306 , n10477 );
    not g21854 ( n654 , n4990 );
    or g21855 ( n25439 , n8422 , n5938 );
    not g21856 ( n486 , n19865 );
    not g21857 ( n21102 , n9669 );
    not g21858 ( n21822 , n15402 );
    and g21859 ( n15333 , n12213 , n10829 );
    not g21860 ( n8333 , n20590 );
    and g21861 ( n26287 , n26363 , n938 );
    or g21862 ( n14312 , n2117 , n19487 );
    not g21863 ( n10749 , n23395 );
    or g21864 ( n10501 , n672 , n2928 );
    not g21865 ( n30535 , n25721 );
    not g21866 ( n2543 , n7358 );
    not g21867 ( n22375 , n18329 );
    xor g21868 ( n4997 , n13605 , n20882 );
    not g21869 ( n3449 , n23965 );
    and g21870 ( n24602 , n17272 , n27759 );
    not g21871 ( n26139 , n12717 );
    not g21872 ( n21115 , n5058 );
    not g21873 ( n9999 , n28927 );
    xnor g21874 ( n2088 , n29362 , n6942 );
    or g21875 ( n21304 , n12174 , n21330 );
    not g21876 ( n5120 , n22042 );
    xnor g21877 ( n16285 , n10155 , n9536 );
    and g21878 ( n25277 , n14350 , n21651 );
    xnor g21879 ( n11372 , n2944 , n15418 );
    or g21880 ( n19782 , n6603 , n3362 );
    or g21881 ( n14009 , n13947 , n15131 );
    not g21882 ( n16042 , n2961 );
    or g21883 ( n4540 , n30887 , n3509 );
    xnor g21884 ( n22185 , n20500 , n26566 );
    or g21885 ( n23426 , n18656 , n12202 );
    nor g21886 ( n18254 , n26106 , n1076 );
    not g21887 ( n27232 , n28031 );
    xnor g21888 ( n17650 , n27615 , n23643 );
    xnor g21889 ( n18877 , n15677 , n3651 );
    not g21890 ( n20862 , n5617 );
    not g21891 ( n7191 , n19484 );
    or g21892 ( n20245 , n27936 , n8510 );
    not g21893 ( n25913 , n31026 );
    nor g21894 ( n18849 , n6681 , n24151 );
    not g21895 ( n18499 , n350 );
    or g21896 ( n3901 , n26564 , n1714 );
    or g21897 ( n16455 , n6914 , n27640 );
    and g21898 ( n29449 , n19411 , n6101 );
    or g21899 ( n28048 , n4821 , n8255 );
    nor g21900 ( n12313 , n11244 , n7670 );
    buf g21901 ( n20967 , n3306 );
    xnor g21902 ( n7076 , n14367 , n13547 );
    xnor g21903 ( n26231 , n12922 , n25695 );
    nor g21904 ( n4600 , n12898 , n7746 );
    and g21905 ( n18552 , n8928 , n13845 );
    not g21906 ( n6613 , n10637 );
    xnor g21907 ( n12018 , n4366 , n17199 );
    xnor g21908 ( n8154 , n24869 , n23167 );
    and g21909 ( n26715 , n2322 , n31395 );
    not g21910 ( n27647 , n23125 );
    not g21911 ( n17084 , n5860 );
    not g21912 ( n23470 , n26115 );
    nor g21913 ( n30117 , n21050 , n26085 );
    xnor g21914 ( n13162 , n8729 , n9130 );
    not g21915 ( n1417 , n22058 );
    nor g21916 ( n1520 , n27448 , n8536 );
    xnor g21917 ( n17415 , n18361 , n1425 );
    xnor g21918 ( n6595 , n31366 , n15436 );
    or g21919 ( n31983 , n11266 , n17721 );
    or g21920 ( n31346 , n17868 , n18056 );
    and g21921 ( n9514 , n8568 , n27932 );
    xnor g21922 ( n6981 , n28790 , n31202 );
    or g21923 ( n9917 , n11085 , n13002 );
    xnor g21924 ( n22504 , n30572 , n29153 );
    not g21925 ( n7409 , n22543 );
    not g21926 ( n24510 , n19300 );
    or g21927 ( n18350 , n1720 , n11082 );
    xnor g21928 ( n7475 , n22673 , n23266 );
    not g21929 ( n20023 , n24439 );
    xnor g21930 ( n5272 , n14263 , n15578 );
    xor g21931 ( n18234 , n10470 , n25190 );
    and g21932 ( n6952 , n28882 , n13665 );
    xnor g21933 ( n26221 , n23535 , n21529 );
    or g21934 ( n31823 , n26523 , n8361 );
    and g21935 ( n910 , n14550 , n4808 );
    and g21936 ( n25238 , n25821 , n23974 );
    and g21937 ( n23790 , n12304 , n32015 );
    nor g21938 ( n25443 , n21185 , n17611 );
    not g21939 ( n10045 , n30579 );
    or g21940 ( n6468 , n21994 , n26268 );
    and g21941 ( n24011 , n19377 , n9433 );
    or g21942 ( n3970 , n4514 , n13026 );
    or g21943 ( n15092 , n22699 , n26634 );
    not g21944 ( n31655 , n21221 );
    xnor g21945 ( n12839 , n5117 , n8792 );
    xnor g21946 ( n18693 , n9940 , n10763 );
    xnor g21947 ( n26408 , n2327 , n31360 );
    xnor g21948 ( n8631 , n27490 , n15060 );
    xnor g21949 ( n31186 , n28774 , n8875 );
    or g21950 ( n22478 , n7909 , n16583 );
    xnor g21951 ( n11245 , n6891 , n6330 );
    xnor g21952 ( n25419 , n31417 , n22139 );
    or g21953 ( n21081 , n22425 , n14986 );
    not g21954 ( n14438 , n8318 );
    and g21955 ( n25342 , n2030 , n30358 );
    nor g21956 ( n12453 , n16347 , n19221 );
    xnor g21957 ( n13116 , n21136 , n18551 );
    xnor g21958 ( n18199 , n5658 , n8197 );
    not g21959 ( n5879 , n18113 );
    xnor g21960 ( n13104 , n13252 , n18851 );
    not g21961 ( n2550 , n1045 );
    xnor g21962 ( n25614 , n11373 , n17981 );
    not g21963 ( n26655 , n8940 );
    or g21964 ( n7196 , n25417 , n874 );
    xnor g21965 ( n21454 , n23038 , n31233 );
    xnor g21966 ( n15760 , n30245 , n11736 );
    xnor g21967 ( n29936 , n4262 , n26114 );
    or g21968 ( n9049 , n30442 , n21657 );
    xnor g21969 ( n19026 , n18756 , n10764 );
    and g21970 ( n21962 , n31537 , n28688 );
    and g21971 ( n21910 , n23238 , n8925 );
    not g21972 ( n11415 , n6153 );
    xnor g21973 ( n7900 , n13474 , n3466 );
    xnor g21974 ( n17281 , n15735 , n18605 );
    not g21975 ( n27133 , n10985 );
    not g21976 ( n17948 , n5912 );
    or g21977 ( n2805 , n6523 , n18971 );
    xnor g21978 ( n11127 , n30143 , n23568 );
    not g21979 ( n13464 , n2925 );
    xnor g21980 ( n5846 , n28409 , n13210 );
    not g21981 ( n12860 , n6783 );
    or g21982 ( n92 , n1866 , n26997 );
    or g21983 ( n12337 , n18193 , n8211 );
    or g21984 ( n15875 , n29933 , n11361 );
    nor g21985 ( n17623 , n16407 , n25711 );
    not g21986 ( n25810 , n18388 );
    and g21987 ( n7397 , n27800 , n7106 );
    or g21988 ( n31003 , n1375 , n7323 );
    not g21989 ( n6916 , n8104 );
    not g21990 ( n18467 , n2340 );
    or g21991 ( n28925 , n10796 , n2600 );
    not g21992 ( n2299 , n26268 );
    and g21993 ( n24880 , n3014 , n15997 );
    not g21994 ( n30761 , n20031 );
    not g21995 ( n19467 , n10514 );
    xnor g21996 ( n11969 , n29437 , n24687 );
    and g21997 ( n28083 , n6170 , n2629 );
    and g21998 ( n7404 , n24738 , n14351 );
    xnor g21999 ( n20888 , n5421 , n12576 );
    and g22000 ( n12494 , n30321 , n18281 );
    or g22001 ( n4336 , n14488 , n23035 );
    xnor g22002 ( n22830 , n13611 , n2081 );
    not g22003 ( n233 , n26192 );
    not g22004 ( n21492 , n24072 );
    nor g22005 ( n22023 , n21506 , n6689 );
    xnor g22006 ( n17028 , n5694 , n28773 );
    not g22007 ( n29541 , n2299 );
    nor g22008 ( n3305 , n9410 , n22499 );
    nor g22009 ( n30449 , n30043 , n29046 );
    or g22010 ( n2602 , n12566 , n196 );
    or g22011 ( n8650 , n30145 , n20368 );
    and g22012 ( n16430 , n2345 , n17465 );
    or g22013 ( n11374 , n18088 , n5865 );
    xnor g22014 ( n1898 , n9939 , n11711 );
    nor g22015 ( n2776 , n9091 , n16740 );
    not g22016 ( n24496 , n3488 );
    nor g22017 ( n15088 , n21979 , n20421 );
    xnor g22018 ( n19162 , n14288 , n2762 );
    or g22019 ( n8072 , n6683 , n10592 );
    not g22020 ( n25493 , n12283 );
    not g22021 ( n8031 , n15845 );
    xnor g22022 ( n18621 , n24625 , n3066 );
    xnor g22023 ( n6532 , n4183 , n4760 );
    not g22024 ( n15242 , n13676 );
    not g22025 ( n6148 , n3828 );
    and g22026 ( n21305 , n20434 , n26258 );
    xnor g22027 ( n1683 , n22499 , n3578 );
    not g22028 ( n26893 , n10873 );
    and g22029 ( n20732 , n17739 , n17109 );
    xnor g22030 ( n23708 , n2434 , n14677 );
    nor g22031 ( n24480 , n15161 , n31648 );
    not g22032 ( n23505 , n4483 );
    or g22033 ( n5667 , n11105 , n18774 );
    nor g22034 ( n1068 , n31755 , n26924 );
    or g22035 ( n28620 , n11785 , n5699 );
    not g22036 ( n21943 , n29966 );
    xnor g22037 ( n28807 , n16541 , n24866 );
    or g22038 ( n3381 , n23786 , n23579 );
    and g22039 ( n25120 , n4816 , n22599 );
    or g22040 ( n3164 , n15491 , n31756 );
    not g22041 ( n31289 , n13363 );
    not g22042 ( n10476 , n3731 );
    and g22043 ( n18766 , n12514 , n2939 );
    xnor g22044 ( n27235 , n22215 , n753 );
    not g22045 ( n23898 , n1720 );
    not g22046 ( n541 , n19521 );
    or g22047 ( n3965 , n9776 , n8987 );
    xnor g22048 ( n3646 , n14919 , n23388 );
    nor g22049 ( n3206 , n26151 , n19396 );
    not g22050 ( n19407 , n10926 );
    or g22051 ( n8204 , n18990 , n6061 );
    or g22052 ( n29074 , n29615 , n31067 );
    or g22053 ( n24434 , n22033 , n17885 );
    not g22054 ( n8732 , n14430 );
    and g22055 ( n2008 , n22937 , n6560 );
    or g22056 ( n16289 , n25079 , n14052 );
    xnor g22057 ( n897 , n27829 , n19255 );
    not g22058 ( n11325 , n30769 );
    or g22059 ( n30512 , n508 , n17645 );
    not g22060 ( n28349 , n2720 );
    or g22061 ( n11029 , n7643 , n1466 );
    and g22062 ( n1435 , n24410 , n4900 );
    xnor g22063 ( n23057 , n10045 , n22422 );
    nor g22064 ( n19475 , n25506 , n1817 );
    xnor g22065 ( n26229 , n6850 , n9824 );
    xnor g22066 ( n18126 , n15577 , n24455 );
    nor g22067 ( n30248 , n28512 , n9378 );
    or g22068 ( n1947 , n12691 , n23295 );
    not g22069 ( n28004 , n11368 );
    not g22070 ( n30374 , n3599 );
    or g22071 ( n8041 , n28584 , n1915 );
    or g22072 ( n19544 , n19405 , n13814 );
    not g22073 ( n5925 , n5863 );
    and g22074 ( n16844 , n8345 , n5066 );
    xnor g22075 ( n15694 , n4674 , n19843 );
    xnor g22076 ( n28220 , n14533 , n3430 );
    or g22077 ( n7739 , n5940 , n11522 );
    not g22078 ( n13057 , n27663 );
    and g22079 ( n25283 , n3437 , n22783 );
    nor g22080 ( n19958 , n27453 , n596 );
    not g22081 ( n2586 , n2174 );
    nor g22082 ( n21626 , n1720 , n21598 );
    and g22083 ( n13026 , n29636 , n31645 );
    or g22084 ( n29922 , n21438 , n8431 );
    not g22085 ( n28428 , n20544 );
    nor g22086 ( n19870 , n3440 , n30095 );
    xnor g22087 ( n18780 , n22340 , n20632 );
    xnor g22088 ( n22920 , n26680 , n18722 );
    or g22089 ( n217 , n20155 , n25347 );
    or g22090 ( n25632 , n853 , n399 );
    or g22091 ( n19969 , n27163 , n4846 );
    not g22092 ( n18092 , n11016 );
    and g22093 ( n13130 , n22508 , n22492 );
    nor g22094 ( n9802 , n27503 , n9445 );
    nor g22095 ( n18967 , n16200 , n7083 );
    not g22096 ( n1179 , n19315 );
    nor g22097 ( n825 , n1346 , n7491 );
    xnor g22098 ( n18853 , n14875 , n28208 );
    xnor g22099 ( n19630 , n5779 , n18307 );
    or g22100 ( n6702 , n30341 , n5743 );
    xor g22101 ( n11434 , n3504 , n12944 );
    xnor g22102 ( n11887 , n29217 , n20311 );
    xnor g22103 ( n31765 , n14450 , n16385 );
    xnor g22104 ( n17821 , n11205 , n9216 );
    nor g22105 ( n18712 , n30121 , n20891 );
    not g22106 ( n18652 , n28428 );
    or g22107 ( n9347 , n26280 , n13810 );
    not g22108 ( n3144 , n13321 );
    not g22109 ( n9652 , n24204 );
    not g22110 ( n12434 , n12075 );
    nor g22111 ( n1788 , n31062 , n11959 );
    xnor g22112 ( n15409 , n11176 , n12158 );
    not g22113 ( n11120 , n26191 );
    xnor g22114 ( n22142 , n18321 , n18400 );
    and g22115 ( n24169 , n22074 , n4646 );
    not g22116 ( n1774 , n12004 );
    nor g22117 ( n16663 , n14954 , n22665 );
    xnor g22118 ( n30659 , n10208 , n22746 );
    and g22119 ( n31704 , n1321 , n18540 );
    or g22120 ( n1927 , n11736 , n9289 );
    or g22121 ( n28550 , n31074 , n4451 );
    or g22122 ( n23149 , n20324 , n18036 );
    or g22123 ( n12997 , n23512 , n4039 );
    and g22124 ( n9444 , n11827 , n12171 );
    not g22125 ( n2985 , n13686 );
    nor g22126 ( n16945 , n25013 , n1350 );
    and g22127 ( n20516 , n16832 , n10751 );
    not g22128 ( n27552 , n19516 );
    nor g22129 ( n2760 , n3753 , n25690 );
    not g22130 ( n28239 , n19846 );
    xnor g22131 ( n15338 , n29658 , n25553 );
    not g22132 ( n3811 , n31543 );
    not g22133 ( n17782 , n26568 );
    or g22134 ( n8502 , n25615 , n19611 );
    or g22135 ( n22117 , n2496 , n11606 );
    and g22136 ( n746 , n6499 , n20124 );
    not g22137 ( n3445 , n20962 );
    not g22138 ( n11032 , n29162 );
    nor g22139 ( n10964 , n22533 , n1316 );
    xnor g22140 ( n20032 , n17307 , n16101 );
    or g22141 ( n8189 , n12627 , n18121 );
    not g22142 ( n20343 , n11073 );
    or g22143 ( n27249 , n17239 , n20217 );
    or g22144 ( n24772 , n14681 , n10252 );
    and g22145 ( n4552 , n28291 , n6336 );
    not g22146 ( n9266 , n31085 );
    not g22147 ( n5988 , n27354 );
    nor g22148 ( n26644 , n5927 , n30146 );
    or g22149 ( n31265 , n27170 , n6288 );
    or g22150 ( n31164 , n17730 , n1120 );
    and g22151 ( n5997 , n3721 , n3250 );
    or g22152 ( n10126 , n7810 , n21962 );
    or g22153 ( n28016 , n5437 , n9637 );
    and g22154 ( n25485 , n30812 , n2250 );
    xnor g22155 ( n23118 , n30602 , n9800 );
    xnor g22156 ( n24479 , n30841 , n20735 );
    xnor g22157 ( n22896 , n2220 , n27389 );
    or g22158 ( n14671 , n22452 , n21952 );
    or g22159 ( n6545 , n11516 , n11089 );
    not g22160 ( n2818 , n23603 );
    not g22161 ( n11283 , n22197 );
    xnor g22162 ( n28674 , n14028 , n31842 );
    xnor g22163 ( n9157 , n11866 , n31783 );
    xnor g22164 ( n6305 , n12934 , n5999 );
    xnor g22165 ( n10657 , n17019 , n12207 );
    not g22166 ( n18767 , n11941 );
    not g22167 ( n30019 , n18905 );
    xnor g22168 ( n19453 , n457 , n14545 );
    not g22169 ( n18328 , n2914 );
    xnor g22170 ( n24901 , n6635 , n106 );
    or g22171 ( n7527 , n20181 , n26529 );
    xnor g22172 ( n14463 , n12643 , n18933 );
    xnor g22173 ( n241 , n22200 , n10737 );
    and g22174 ( n24542 , n10510 , n7840 );
    xnor g22175 ( n5484 , n11308 , n27708 );
    and g22176 ( n7165 , n4741 , n31063 );
    or g22177 ( n18805 , n1653 , n11441 );
    not g22178 ( n10463 , n31313 );
    not g22179 ( n3115 , n7645 );
    not g22180 ( n28368 , n28535 );
    not g22181 ( n21607 , n22075 );
    not g22182 ( n21901 , n9566 );
    not g22183 ( n17966 , n32020 );
    or g22184 ( n1398 , n29106 , n4886 );
    nor g22185 ( n11897 , n3004 , n22493 );
    or g22186 ( n26427 , n18080 , n7725 );
    nor g22187 ( n31583 , n12205 , n11607 );
    and g22188 ( n1832 , n15475 , n22096 );
    or g22189 ( n24749 , n10446 , n31994 );
    nor g22190 ( n20675 , n27322 , n9455 );
    or g22191 ( n24706 , n30210 , n19048 );
    xnor g22192 ( n4993 , n6392 , n21290 );
    xnor g22193 ( n31150 , n27318 , n1404 );
    not g22194 ( n26991 , n12468 );
    or g22195 ( n27931 , n13169 , n1595 );
    not g22196 ( n18412 , n20486 );
    not g22197 ( n406 , n23372 );
    or g22198 ( n21193 , n31940 , n24953 );
    not g22199 ( n23699 , n16264 );
    xor g22200 ( n21855 , n4289 , n11255 );
    xnor g22201 ( n25848 , n30908 , n7692 );
    or g22202 ( n25762 , n22947 , n26666 );
    or g22203 ( n11422 , n20190 , n20404 );
    and g22204 ( n25612 , n8389 , n25021 );
    xnor g22205 ( n11945 , n1177 , n1692 );
    not g22206 ( n9121 , n18691 );
    xnor g22207 ( n21718 , n31806 , n26598 );
    not g22208 ( n28390 , n16649 );
    or g22209 ( n8237 , n11776 , n16153 );
    and g22210 ( n7522 , n3692 , n12920 );
    xnor g22211 ( n3417 , n25351 , n28375 );
    and g22212 ( n22811 , n4389 , n23837 );
    not g22213 ( n5485 , n20130 );
    and g22214 ( n6173 , n29468 , n17290 );
    nor g22215 ( n511 , n21030 , n4432 );
    xor g22216 ( n3661 , n28585 , n7849 );
    buf g22217 ( n16083 , n5820 );
    and g22218 ( n9728 , n30086 , n28817 );
    and g22219 ( n25478 , n23060 , n25972 );
    and g22220 ( n15562 , n7233 , n27781 );
    or g22221 ( n23501 , n16571 , n7595 );
    and g22222 ( n28505 , n25217 , n3375 );
    xnor g22223 ( n12577 , n20942 , n1591 );
    not g22224 ( n1050 , n18296 );
    not g22225 ( n18216 , n26082 );
    xnor g22226 ( n19153 , n30287 , n16113 );
    xnor g22227 ( n5666 , n30678 , n11169 );
    xnor g22228 ( n28572 , n6798 , n30238 );
    xnor g22229 ( n20895 , n8038 , n9610 );
    xnor g22230 ( n4195 , n25611 , n17504 );
    not g22231 ( n7603 , n11513 );
    not g22232 ( n1624 , n6559 );
    or g22233 ( n31157 , n4517 , n24865 );
    and g22234 ( n1714 , n1402 , n271 );
    or g22235 ( n5110 , n28904 , n25281 );
    xnor g22236 ( n10529 , n10633 , n2447 );
    xnor g22237 ( n729 , n25286 , n24786 );
    not g22238 ( n16029 , n6139 );
    not g22239 ( n10960 , n13065 );
    or g22240 ( n31235 , n30822 , n26298 );
    nor g22241 ( n10449 , n30434 , n20104 );
    not g22242 ( n29873 , n24197 );
    not g22243 ( n1032 , n6141 );
    not g22244 ( n14314 , n13864 );
    xor g22245 ( n16845 , n17569 , n28675 );
    or g22246 ( n13098 , n25486 , n8463 );
    not g22247 ( n22072 , n24965 );
    xnor g22248 ( n22702 , n14650 , n374 );
    or g22249 ( n26719 , n18951 , n9086 );
    and g22250 ( n4231 , n18786 , n25732 );
    or g22251 ( n16966 , n15755 , n19368 );
    xnor g22252 ( n17885 , n22770 , n4709 );
    or g22253 ( n21900 , n13901 , n26903 );
    and g22254 ( n25148 , n23004 , n3354 );
    xnor g22255 ( n21997 , n15268 , n16347 );
    xnor g22256 ( n28096 , n975 , n1709 );
    or g22257 ( n23913 , n5430 , n23454 );
    xnor g22258 ( n27442 , n20986 , n9806 );
    not g22259 ( n10194 , n19572 );
    not g22260 ( n10029 , n1131 );
    and g22261 ( n16353 , n24347 , n9958 );
    xnor g22262 ( n27214 , n29184 , n19529 );
    not g22263 ( n11674 , n2963 );
    and g22264 ( n19966 , n29231 , n8833 );
    not g22265 ( n21764 , n31450 );
    xnor g22266 ( n9842 , n3871 , n17749 );
    and g22267 ( n11207 , n4438 , n15099 );
    or g22268 ( n23370 , n3295 , n23541 );
    nor g22269 ( n6317 , n26799 , n11052 );
    nor g22270 ( n7791 , n11729 , n568 );
    or g22271 ( n30175 , n12409 , n16331 );
    xnor g22272 ( n5080 , n20774 , n28009 );
    xnor g22273 ( n2676 , n2808 , n22549 );
    or g22274 ( n25754 , n20732 , n14031 );
    or g22275 ( n30462 , n20445 , n13804 );
    or g22276 ( n19234 , n346 , n20382 );
    or g22277 ( n15741 , n7001 , n17494 );
    xnor g22278 ( n31540 , n18606 , n27832 );
    not g22279 ( n14724 , n25758 );
    xnor g22280 ( n29502 , n3858 , n20116 );
    and g22281 ( n13558 , n10316 , n8781 );
    and g22282 ( n21518 , n12263 , n3997 );
    or g22283 ( n28285 , n14176 , n6860 );
    not g22284 ( n23671 , n15514 );
    xnor g22285 ( n19202 , n13341 , n22896 );
    or g22286 ( n16752 , n12749 , n1929 );
    not g22287 ( n12756 , n4414 );
    not g22288 ( n21778 , n18619 );
    xnor g22289 ( n17818 , n24989 , n21312 );
    nor g22290 ( n19753 , n8348 , n15714 );
    not g22291 ( n26073 , n31092 );
    or g22292 ( n15121 , n10574 , n5257 );
    xnor g22293 ( n2851 , n6566 , n530 );
    not g22294 ( n10364 , n20769 );
    or g22295 ( n24401 , n13515 , n10181 );
    nor g22296 ( n7784 , n2447 , n10633 );
    nor g22297 ( n13671 , n5573 , n5528 );
    not g22298 ( n21401 , n28141 );
    not g22299 ( n3375 , n27416 );
    or g22300 ( n1249 , n13229 , n1581 );
    not g22301 ( n1102 , n15493 );
    or g22302 ( n27890 , n8097 , n6866 );
    xnor g22303 ( n25742 , n14570 , n9906 );
    or g22304 ( n1295 , n8133 , n30276 );
    xnor g22305 ( n4702 , n15758 , n13833 );
    xnor g22306 ( n17833 , n3170 , n13833 );
    or g22307 ( n13452 , n1177 , n6416 );
    and g22308 ( n497 , n30308 , n19363 );
    and g22309 ( n32017 , n10849 , n17451 );
    nor g22310 ( n30441 , n23255 , n7439 );
    not g22311 ( n13555 , n29785 );
    xnor g22312 ( n18648 , n2963 , n22233 );
    or g22313 ( n16798 , n26628 , n16908 );
    xnor g22314 ( n24360 , n26635 , n23081 );
    and g22315 ( n27756 , n5613 , n18912 );
    not g22316 ( n20508 , n23330 );
    xnor g22317 ( n29348 , n15587 , n24037 );
    not g22318 ( n25194 , n29083 );
    or g22319 ( n11040 , n10434 , n32005 );
    and g22320 ( n16929 , n22200 , n10737 );
    and g22321 ( n17566 , n29775 , n8511 );
    not g22322 ( n5664 , n30524 );
    xnor g22323 ( n18504 , n7223 , n18582 );
    not g22324 ( n4523 , n16963 );
    or g22325 ( n4912 , n9861 , n29543 );
    or g22326 ( n20333 , n26241 , n26453 );
    xnor g22327 ( n29976 , n8522 , n24113 );
    and g22328 ( n7883 , n20558 , n6896 );
    not g22329 ( n17455 , n3307 );
    and g22330 ( n10426 , n2942 , n26161 );
    and g22331 ( n13626 , n22869 , n13851 );
    not g22332 ( n30209 , n11724 );
    nor g22333 ( n20070 , n18203 , n17813 );
    nor g22334 ( n7311 , n14670 , n14962 );
    xnor g22335 ( n12679 , n20870 , n4350 );
    xnor g22336 ( n18675 , n19705 , n16088 );
    nor g22337 ( n18862 , n28006 , n3454 );
    xnor g22338 ( n19607 , n11256 , n1088 );
    and g22339 ( n24253 , n25465 , n5595 );
    and g22340 ( n11759 , n12771 , n5149 );
    and g22341 ( n10512 , n19470 , n9471 );
    and g22342 ( n16668 , n31870 , n8304 );
    not g22343 ( n965 , n10433 );
    nor g22344 ( n19392 , n17302 , n9829 );
    xnor g22345 ( n23382 , n29056 , n20736 );
    xnor g22346 ( n18037 , n31860 , n235 );
    not g22347 ( n23980 , n5963 );
    xnor g22348 ( n4317 , n29724 , n19144 );
    xnor g22349 ( n3981 , n23537 , n4887 );
    not g22350 ( n8172 , n24824 );
    not g22351 ( n15172 , n25585 );
    or g22352 ( n17972 , n14111 , n31054 );
    not g22353 ( n23547 , n4780 );
    not g22354 ( n4258 , n28523 );
    and g22355 ( n4837 , n10026 , n22436 );
    not g22356 ( n24935 , n27789 );
    not g22357 ( n22942 , n2333 );
    xnor g22358 ( n22607 , n12806 , n13514 );
    not g22359 ( n17006 , n15772 );
    not g22360 ( n3582 , n1857 );
    not g22361 ( n13749 , n11912 );
    xnor g22362 ( n15260 , n29245 , n5150 );
    not g22363 ( n5659 , n14869 );
    nor g22364 ( n18102 , n19554 , n29482 );
    not g22365 ( n6943 , n29550 );
    nor g22366 ( n2576 , n11851 , n25344 );
    not g22367 ( n28962 , n28983 );
    nor g22368 ( n14046 , n3611 , n2918 );
    or g22369 ( n19191 , n6732 , n28819 );
    xor g22370 ( n12028 , n14340 , n10393 );
    not g22371 ( n29296 , n5166 );
    and g22372 ( n7292 , n17769 , n10052 );
    or g22373 ( n23888 , n18378 , n18070 );
    not g22374 ( n16128 , n22875 );
    or g22375 ( n3405 , n29974 , n27867 );
    or g22376 ( n3337 , n12933 , n5489 );
    not g22377 ( n13582 , n18208 );
    and g22378 ( n4869 , n12459 , n12645 );
    or g22379 ( n1369 , n3059 , n9066 );
    nor g22380 ( n13994 , n30171 , n7732 );
    xnor g22381 ( n16204 , n10954 , n23597 );
    not g22382 ( n22033 , n31028 );
    not g22383 ( n18889 , n6543 );
    or g22384 ( n20838 , n2511 , n15584 );
    and g22385 ( n3927 , n25316 , n28812 );
    xnor g22386 ( n7548 , n3684 , n26012 );
    and g22387 ( n28653 , n22210 , n14106 );
    and g22388 ( n11767 , n25434 , n7084 );
    and g22389 ( n28182 , n19677 , n501 );
    nor g22390 ( n27760 , n20181 , n25188 );
    xnor g22391 ( n9806 , n29094 , n2404 );
    or g22392 ( n613 , n25793 , n2665 );
    not g22393 ( n15970 , n11583 );
    or g22394 ( n1047 , n2643 , n12808 );
    nor g22395 ( n23512 , n13751 , n15382 );
    xnor g22396 ( n12766 , n27539 , n4160 );
    and g22397 ( n6496 , n4549 , n5764 );
    xnor g22398 ( n5083 , n385 , n17660 );
    xnor g22399 ( n8126 , n14882 , n27064 );
    not g22400 ( n19463 , n28942 );
    xnor g22401 ( n6827 , n3053 , n27407 );
    or g22402 ( n11451 , n29177 , n23237 );
    xnor g22403 ( n13102 , n10219 , n12488 );
    and g22404 ( n15524 , n722 , n12314 );
    or g22405 ( n11442 , n22611 , n5810 );
    and g22406 ( n14614 , n17629 , n30224 );
    or g22407 ( n30241 , n3182 , n6305 );
    or g22408 ( n714 , n95 , n19070 );
    not g22409 ( n28346 , n19344 );
    xnor g22410 ( n14939 , n10390 , n29986 );
    or g22411 ( n1885 , n29841 , n29951 );
    xnor g22412 ( n13154 , n21174 , n5345 );
    nor g22413 ( n19908 , n3080 , n11706 );
    xnor g22414 ( n6350 , n24507 , n18718 );
    xnor g22415 ( n17864 , n632 , n12364 );
    not g22416 ( n23480 , n30793 );
    or g22417 ( n3982 , n4014 , n7789 );
    not g22418 ( n25033 , n18373 );
    nor g22419 ( n7035 , n7055 , n23365 );
    or g22420 ( n14247 , n20986 , n4715 );
    not g22421 ( n14097 , n27954 );
    not g22422 ( n14415 , n12705 );
    or g22423 ( n6353 , n30848 , n13694 );
    or g22424 ( n24346 , n29949 , n8574 );
    not g22425 ( n19345 , n21107 );
    and g22426 ( n14061 , n14619 , n16574 );
    not g22427 ( n223 , n21891 );
    and g22428 ( n5577 , n14654 , n15051 );
    and g22429 ( n6755 , n4765 , n28147 );
    buf g22430 ( n23184 , n21588 );
    and g22431 ( n23686 , n29461 , n1611 );
    not g22432 ( n5115 , n6014 );
    and g22433 ( n2817 , n9422 , n11456 );
    and g22434 ( n26930 , n25694 , n28838 );
    not g22435 ( n24766 , n11284 );
    or g22436 ( n19967 , n9306 , n25912 );
    buf g22437 ( n18612 , n24072 );
    nor g22438 ( n20352 , n11736 , n22043 );
    and g22439 ( n17931 , n31022 , n10360 );
    or g22440 ( n25105 , n9479 , n2328 );
    nor g22441 ( n15394 , n10960 , n5498 );
    not g22442 ( n23992 , n5896 );
    and g22443 ( n22571 , n5031 , n3533 );
    not g22444 ( n27491 , n16406 );
    xnor g22445 ( n10159 , n24280 , n2200 );
    or g22446 ( n216 , n29561 , n30880 );
    and g22447 ( n15248 , n5761 , n19442 );
    or g22448 ( n11350 , n29771 , n17096 );
    not g22449 ( n3420 , n835 );
    xnor g22450 ( n9568 , n406 , n15798 );
    xnor g22451 ( n24251 , n25793 , n2665 );
    not g22452 ( n16149 , n17900 );
    or g22453 ( n8372 , n13296 , n13666 );
    xnor g22454 ( n14998 , n1418 , n4372 );
    and g22455 ( n31476 , n4410 , n24794 );
    not g22456 ( n27729 , n16291 );
    not g22457 ( n514 , n22568 );
    not g22458 ( n3824 , n1798 );
    not g22459 ( n31271 , n3029 );
    not g22460 ( n316 , n31631 );
    not g22461 ( n18881 , n18850 );
    not g22462 ( n12451 , n17896 );
    xnor g22463 ( n5027 , n10007 , n7299 );
    or g22464 ( n26994 , n14227 , n13526 );
    and g22465 ( n12506 , n9667 , n19060 );
    not g22466 ( n14955 , n19408 );
    xnor g22467 ( n30310 , n18579 , n4292 );
    not g22468 ( n21947 , n23410 );
    and g22469 ( n17965 , n7251 , n5815 );
    xnor g22470 ( n20196 , n25093 , n2301 );
    and g22471 ( n22499 , n17412 , n15647 );
    and g22472 ( n11196 , n29181 , n23021 );
    and g22473 ( n8444 , n12917 , n18290 );
    or g22474 ( n31052 , n3765 , n12879 );
    not g22475 ( n12233 , n22777 );
    xnor g22476 ( n9632 , n31195 , n15779 );
    or g22477 ( n26749 , n10114 , n3782 );
    and g22478 ( n27861 , n18523 , n4331 );
    xnor g22479 ( n8497 , n23218 , n19538 );
    not g22480 ( n17912 , n11010 );
    buf g22481 ( n30574 , n31386 );
    nor g22482 ( n24657 , n5561 , n1067 );
    xnor g22483 ( n2978 , n1551 , n5299 );
    nor g22484 ( n11446 , n2483 , n5384 );
    or g22485 ( n6357 , n22512 , n23369 );
    nor g22486 ( n26922 , n2588 , n6107 );
    or g22487 ( n29809 , n2213 , n25117 );
    not g22488 ( n8571 , n28637 );
    and g22489 ( n14402 , n8635 , n30802 );
    xnor g22490 ( n30472 , n26533 , n30498 );
    xnor g22491 ( n26848 , n26996 , n11065 );
    or g22492 ( n12301 , n9287 , n24326 );
    xnor g22493 ( n15050 , n21947 , n2072 );
    and g22494 ( n14525 , n3593 , n5826 );
    xnor g22495 ( n15995 , n11149 , n4055 );
    not g22496 ( n2777 , n19599 );
    or g22497 ( n31322 , n16521 , n23640 );
    or g22498 ( n27815 , n14690 , n17037 );
    not g22499 ( n12373 , n15219 );
    xnor g22500 ( n15580 , n2747 , n28821 );
    and g22501 ( n27633 , n4301 , n17409 );
    not g22502 ( n28524 , n18065 );
    and g22503 ( n24994 , n5956 , n30072 );
    not g22504 ( n2914 , n25393 );
    not g22505 ( n5361 , n15558 );
    not g22506 ( n16444 , n2855 );
    nor g22507 ( n6434 , n84 , n6803 );
    xnor g22508 ( n8378 , n22384 , n16549 );
    and g22509 ( n5285 , n12432 , n15605 );
    and g22510 ( n13878 , n15023 , n10586 );
    not g22511 ( n2965 , n26324 );
    or g22512 ( n30125 , n13678 , n5552 );
    xnor g22513 ( n28336 , n17341 , n14175 );
    or g22514 ( n30644 , n3554 , n10307 );
    xnor g22515 ( n21584 , n21918 , n21771 );
    or g22516 ( n2900 , n22219 , n3718 );
    and g22517 ( n25459 , n22588 , n9953 );
    xnor g22518 ( n31037 , n16276 , n17286 );
    or g22519 ( n13806 , n2960 , n2553 );
    not g22520 ( n28721 , n28795 );
    and g22521 ( n4138 , n29059 , n24184 );
    or g22522 ( n8979 , n30895 , n26341 );
    xnor g22523 ( n20246 , n17728 , n12255 );
    not g22524 ( n16508 , n14503 );
    or g22525 ( n20300 , n19274 , n5868 );
    nor g22526 ( n9123 , n7209 , n27591 );
    nor g22527 ( n25074 , n24153 , n12188 );
    and g22528 ( n22131 , n12096 , n16193 );
    nor g22529 ( n9930 , n31108 , n20765 );
    or g22530 ( n15011 , n14513 , n19790 );
    not g22531 ( n15101 , n6532 );
    xnor g22532 ( n7225 , n29275 , n31751 );
    or g22533 ( n10248 , n1736 , n15272 );
    not g22534 ( n25702 , n14195 );
    and g22535 ( n1446 , n9562 , n2168 );
    and g22536 ( n31533 , n4444 , n2039 );
    and g22537 ( n4354 , n17091 , n30222 );
    nor g22538 ( n10675 , n2124 , n9838 );
    and g22539 ( n9501 , n29381 , n9893 );
    xnor g22540 ( n31590 , n6041 , n12816 );
    not g22541 ( n12154 , n10054 );
    nor g22542 ( n11728 , n24775 , n12979 );
    or g22543 ( n30551 , n15784 , n21884 );
    or g22544 ( n9076 , n30458 , n8622 );
    and g22545 ( n25903 , n2464 , n28409 );
    not g22546 ( n17895 , n30124 );
    and g22547 ( n15456 , n26962 , n11115 );
    xnor g22548 ( n18613 , n26082 , n23342 );
    nor g22549 ( n16895 , n12105 , n16322 );
    or g22550 ( n18414 , n16609 , n2176 );
    or g22551 ( n19249 , n6355 , n1475 );
    nor g22552 ( n4232 , n26358 , n20644 );
    xnor g22553 ( n3686 , n19789 , n17818 );
    xnor g22554 ( n3946 , n12970 , n14477 );
    and g22555 ( n1430 , n31001 , n629 );
    or g22556 ( n15139 , n8943 , n14938 );
    not g22557 ( n28575 , n24819 );
    not g22558 ( n7357 , n26670 );
    or g22559 ( n31991 , n11990 , n28095 );
    or g22560 ( n29067 , n18667 , n23817 );
    xnor g22561 ( n13257 , n1526 , n5834 );
    xnor g22562 ( n26624 , n17925 , n6345 );
    and g22563 ( n6522 , n30317 , n27664 );
    nor g22564 ( n17736 , n12713 , n2668 );
    buf g22565 ( n24584 , n8478 );
    not g22566 ( n17079 , n12192 );
    or g22567 ( n26681 , n8768 , n19128 );
    and g22568 ( n23383 , n21503 , n971 );
    xnor g22569 ( n17464 , n17302 , n28180 );
    and g22570 ( n3703 , n13856 , n10584 );
    nor g22571 ( n24218 , n30664 , n17842 );
    or g22572 ( n25327 , n3080 , n9591 );
    not g22573 ( n1078 , n11462 );
    and g22574 ( n3116 , n25041 , n9003 );
    or g22575 ( n4985 , n29837 , n31110 );
    not g22576 ( n30253 , n15092 );
    nor g22577 ( n7970 , n6069 , n28524 );
    or g22578 ( n2884 , n6146 , n27816 );
    or g22579 ( n6668 , n31743 , n16145 );
    not g22580 ( n13197 , n28333 );
    xnor g22581 ( n15360 , n2186 , n3791 );
    or g22582 ( n30615 , n21753 , n13461 );
    not g22583 ( n26805 , n19896 );
    and g22584 ( n7173 , n21762 , n186 );
    xor g22585 ( n24612 , n24174 , n953 );
    or g22586 ( n17817 , n54 , n1777 );
    and g22587 ( n3353 , n17937 , n25975 );
    nor g22588 ( n19285 , n17220 , n20178 );
    xnor g22589 ( n11470 , n26633 , n13700 );
    or g22590 ( n21827 , n32019 , n7420 );
    not g22591 ( n23024 , n21322 );
    xnor g22592 ( n19921 , n3367 , n11984 );
    nor g22593 ( n29498 , n3488 , n13888 );
    not g22594 ( n27435 , n29949 );
    not g22595 ( n25472 , n4915 );
    and g22596 ( n5163 , n1916 , n2083 );
    xnor g22597 ( n21290 , n15641 , n30909 );
    xnor g22598 ( n13060 , n9068 , n13222 );
    or g22599 ( n20658 , n4090 , n1408 );
    or g22600 ( n25081 , n24783 , n25011 );
    xnor g22601 ( n5052 , n27992 , n21192 );
    not g22602 ( n19427 , n23052 );
    not g22603 ( n20828 , n25306 );
    xnor g22604 ( n28603 , n2928 , n28518 );
    not g22605 ( n29125 , n32011 );
    xnor g22606 ( n22574 , n29271 , n6144 );
    or g22607 ( n25622 , n11247 , n5262 );
    xnor g22608 ( n29553 , n13014 , n3369 );
    not g22609 ( n17205 , n2358 );
    nor g22610 ( n30716 , n16108 , n27581 );
    not g22611 ( n24336 , n15813 );
    not g22612 ( n27899 , n12364 );
    xnor g22613 ( n6471 , n14103 , n31171 );
    xnor g22614 ( n1977 , n4512 , n19092 );
    not g22615 ( n13433 , n3142 );
    or g22616 ( n2979 , n10609 , n29788 );
    not g22617 ( n3065 , n8157 );
    or g22618 ( n1076 , n5687 , n15430 );
    and g22619 ( n29013 , n24370 , n23586 );
    xnor g22620 ( n20075 , n23868 , n20788 );
    or g22621 ( n24868 , n4430 , n7142 );
    and g22622 ( n12723 , n21745 , n13997 );
    or g22623 ( n21471 , n22461 , n2868 );
    xnor g22624 ( n25690 , n26215 , n15482 );
    and g22625 ( n12505 , n1662 , n14043 );
    or g22626 ( n4753 , n13604 , n25072 );
    not g22627 ( n6086 , n4408 );
    not g22628 ( n4330 , n6305 );
    and g22629 ( n14963 , n9143 , n9308 );
    xnor g22630 ( n19358 , n21627 , n18769 );
    xnor g22631 ( n10797 , n12084 , n22294 );
    not g22632 ( n18538 , n23185 );
    and g22633 ( n22215 , n17450 , n7388 );
    and g22634 ( n21000 , n854 , n29378 );
    not g22635 ( n30594 , n27126 );
    xnor g22636 ( n26430 , n6535 , n10860 );
    not g22637 ( n11322 , n24161 );
    or g22638 ( n22700 , n12309 , n13580 );
    or g22639 ( n1136 , n9265 , n19367 );
    or g22640 ( n71 , n19637 , n26347 );
    or g22641 ( n23215 , n19025 , n12988 );
    or g22642 ( n18628 , n24171 , n21631 );
    or g22643 ( n146 , n19443 , n29150 );
    or g22644 ( n26421 , n17191 , n16820 );
    not g22645 ( n16716 , n15334 );
    nor g22646 ( n1737 , n2898 , n17305 );
    not g22647 ( n2553 , n30161 );
    or g22648 ( n25775 , n4325 , n8678 );
    not g22649 ( n24863 , n13184 );
    or g22650 ( n30493 , n28431 , n31156 );
    or g22651 ( n21109 , n1014 , n6348 );
    and g22652 ( n31610 , n1294 , n20299 );
    not g22653 ( n17667 , n28593 );
    or g22654 ( n5855 , n4545 , n29625 );
    xnor g22655 ( n21530 , n28247 , n21122 );
    or g22656 ( n2412 , n16998 , n13660 );
    not g22657 ( n28489 , n12233 );
    nor g22658 ( n18568 , n2963 , n1913 );
    or g22659 ( n2096 , n19066 , n25675 );
    xnor g22660 ( n15895 , n31865 , n12645 );
    xnor g22661 ( n13958 , n22906 , n26459 );
    not g22662 ( n24265 , n9174 );
    and g22663 ( n12209 , n2845 , n14926 );
    xnor g22664 ( n28386 , n16933 , n24266 );
    nor g22665 ( n20292 , n25046 , n31759 );
    or g22666 ( n25107 , n8336 , n17002 );
    not g22667 ( n31333 , n1671 );
    nor g22668 ( n8950 , n24387 , n11552 );
    nor g22669 ( n4519 , n2001 , n8610 );
    not g22670 ( n21690 , n14901 );
    and g22671 ( n12811 , n5918 , n27542 );
    or g22672 ( n4309 , n427 , n8046 );
    and g22673 ( n31506 , n28308 , n17401 );
    not g22674 ( n31394 , n9472 );
    or g22675 ( n25015 , n23383 , n3168 );
    nor g22676 ( n24745 , n8584 , n28962 );
    xnor g22677 ( n5737 , n19116 , n1818 );
    not g22678 ( n7395 , n31982 );
    or g22679 ( n3468 , n31338 , n12468 );
    xnor g22680 ( n24182 , n24266 , n14324 );
    not g22681 ( n7042 , n19839 );
    and g22682 ( n23454 , n21985 , n30628 );
    or g22683 ( n24928 , n4791 , n7838 );
    or g22684 ( n13816 , n31952 , n28059 );
    xnor g22685 ( n6895 , n17029 , n547 );
    xnor g22686 ( n17233 , n18218 , n14851 );
    not g22687 ( n4551 , n20215 );
    and g22688 ( n24300 , n27100 , n9452 );
    xnor g22689 ( n23111 , n22003 , n31199 );
    xnor g22690 ( n8875 , n20112 , n26858 );
    or g22691 ( n25845 , n6614 , n27404 );
    not g22692 ( n12198 , n9935 );
    not g22693 ( n20820 , n3010 );
    nor g22694 ( n30473 , n26306 , n7611 );
    and g22695 ( n21992 , n29729 , n18032 );
    xnor g22696 ( n7808 , n20973 , n16677 );
    xnor g22697 ( n14479 , n9056 , n14003 );
    or g22698 ( n21283 , n3087 , n21367 );
    xnor g22699 ( n18660 , n9327 , n25820 );
    or g22700 ( n22457 , n13403 , n20711 );
    xnor g22701 ( n2373 , n3064 , n11519 );
    xnor g22702 ( n18590 , n23190 , n1677 );
    not g22703 ( n5332 , n29641 );
    or g22704 ( n24668 , n21488 , n15078 );
    and g22705 ( n12371 , n24570 , n8245 );
    xnor g22706 ( n4052 , n29823 , n11 );
    or g22707 ( n26175 , n12423 , n8932 );
    not g22708 ( n19375 , n19557 );
    not g22709 ( n27389 , n23069 );
    and g22710 ( n645 , n22654 , n16230 );
    nor g22711 ( n27073 , n11226 , n27693 );
    and g22712 ( n173 , n26279 , n26957 );
    xnor g22713 ( n8927 , n5613 , n14105 );
    and g22714 ( n6284 , n21618 , n13327 );
    xnor g22715 ( n24916 , n6814 , n3665 );
    not g22716 ( n22654 , n7450 );
    or g22717 ( n12731 , n3386 , n16517 );
    xor g22718 ( n30974 , n30894 , n25535 );
    nor g22719 ( n11855 , n12318 , n11481 );
    xnor g22720 ( n25214 , n15080 , n3780 );
    and g22721 ( n4303 , n13775 , n31177 );
    xor g22722 ( n5451 , n10591 , n27497 );
    or g22723 ( n19800 , n13883 , n29957 );
    or g22724 ( n25090 , n14636 , n24784 );
    not g22725 ( n31600 , n30987 );
    or g22726 ( n24808 , n31589 , n2718 );
    or g22727 ( n19020 , n22939 , n6617 );
    or g22728 ( n2045 , n2910 , n21600 );
    xnor g22729 ( n3489 , n20632 , n28634 );
    xnor g22730 ( n3593 , n27038 , n11550 );
    xnor g22731 ( n2055 , n14962 , n11060 );
    not g22732 ( n23842 , n12399 );
    xnor g22733 ( n7492 , n2844 , n21132 );
    nor g22734 ( n356 , n24615 , n10880 );
    and g22735 ( n13166 , n28151 , n11605 );
    and g22736 ( n8675 , n25984 , n27537 );
    or g22737 ( n29211 , n15015 , n24705 );
    xnor g22738 ( n5273 , n12510 , n29734 );
    or g22739 ( n16868 , n26032 , n18258 );
    not g22740 ( n4274 , n7705 );
    xnor g22741 ( n8054 , n28093 , n13781 );
    xnor g22742 ( n25984 , n24543 , n21445 );
    xnor g22743 ( n29427 , n16320 , n4829 );
    not g22744 ( n8529 , n862 );
    and g22745 ( n28072 , n437 , n26178 );
    and g22746 ( n27738 , n29738 , n21167 );
    or g22747 ( n17538 , n12882 , n30254 );
    xnor g22748 ( n18637 , n26974 , n2001 );
    or g22749 ( n3575 , n19300 , n11624 );
    xnor g22750 ( n26885 , n22480 , n31278 );
    or g22751 ( n18563 , n28946 , n2476 );
    not g22752 ( n22355 , n24185 );
    or g22753 ( n23331 , n2782 , n22775 );
    or g22754 ( n22394 , n16391 , n10718 );
    and g22755 ( n9107 , n28015 , n6991 );
    or g22756 ( n11208 , n20723 , n2102 );
    and g22757 ( n24823 , n4211 , n4758 );
    and g22758 ( n23390 , n21153 , n15500 );
    not g22759 ( n12550 , n6626 );
    not g22760 ( n7051 , n29878 );
    or g22761 ( n19817 , n8879 , n1510 );
    or g22762 ( n638 , n18287 , n7537 );
    not g22763 ( n11645 , n6874 );
    nor g22764 ( n30677 , n7552 , n30939 );
    not g22765 ( n15245 , n5459 );
    xnor g22766 ( n11609 , n16856 , n154 );
    xor g22767 ( n6322 , n20302 , n28029 );
    or g22768 ( n30192 , n6708 , n7820 );
    buf g22769 ( n24369 , n9490 );
    xnor g22770 ( n16584 , n25056 , n6750 );
    or g22771 ( n10987 , n18033 , n1582 );
    xnor g22772 ( n22541 , n22435 , n29398 );
    xnor g22773 ( n12681 , n30581 , n29208 );
    not g22774 ( n21002 , n15588 );
    not g22775 ( n22234 , n31910 );
    not g22776 ( n11435 , n14067 );
    xnor g22777 ( n31332 , n2449 , n28510 );
    or g22778 ( n20551 , n5908 , n22052 );
    xnor g22779 ( n6543 , n2121 , n8920 );
    or g22780 ( n13198 , n18739 , n21163 );
    and g22781 ( n27606 , n12507 , n23762 );
    not g22782 ( n13977 , n3719 );
    or g22783 ( n17410 , n10656 , n14674 );
    xnor g22784 ( n21814 , n19171 , n7009 );
    or g22785 ( n26134 , n29359 , n25554 );
    not g22786 ( n24268 , n21741 );
    xnor g22787 ( n30370 , n26364 , n9655 );
    not g22788 ( n13993 , n7662 );
    and g22789 ( n698 , n29357 , n621 );
    nor g22790 ( n4957 , n21629 , n30301 );
    and g22791 ( n18592 , n10745 , n9027 );
    or g22792 ( n27191 , n18776 , n7039 );
    nor g22793 ( n8677 , n13275 , n23756 );
    xnor g22794 ( n17133 , n15635 , n29132 );
    and g22795 ( n5959 , n22774 , n1724 );
    not g22796 ( n31935 , n13375 );
    or g22797 ( n4866 , n17600 , n6587 );
    not g22798 ( n3884 , n17479 );
    and g22799 ( n4874 , n24466 , n25703 );
    or g22800 ( n12044 , n17856 , n23432 );
    xnor g22801 ( n9490 , n25440 , n19306 );
    and g22802 ( n29027 , n25619 , n20619 );
    or g22803 ( n28586 , n19108 , n2228 );
    or g22804 ( n5548 , n9176 , n26902 );
    not g22805 ( n28794 , n4168 );
    nor g22806 ( n31403 , n9239 , n14328 );
    and g22807 ( n20711 , n20609 , n12257 );
    or g22808 ( n22638 , n19540 , n15851 );
    nor g22809 ( n332 , n26961 , n942 );
    nor g22810 ( n4394 , n22867 , n16920 );
    nor g22811 ( n13180 , n17478 , n18310 );
    and g22812 ( n20873 , n12648 , n1103 );
    not g22813 ( n12941 , n29261 );
    or g22814 ( n25224 , n580 , n4523 );
    and g22815 ( n21011 , n11213 , n9573 );
    or g22816 ( n5206 , n9935 , n679 );
    not g22817 ( n10844 , n1381 );
    not g22818 ( n3505 , n14887 );
    xor g22819 ( n28643 , n31355 , n13859 );
    not g22820 ( n16806 , n27733 );
    or g22821 ( n18580 , n21301 , n15208 );
    xnor g22822 ( n11531 , n15315 , n8988 );
    or g22823 ( n8339 , n5042 , n3881 );
    not g22824 ( n2432 , n26700 );
    or g22825 ( n11460 , n17845 , n28093 );
    or g22826 ( n22061 , n3681 , n2929 );
    xnor g22827 ( n28116 , n9007 , n3229 );
    not g22828 ( n24445 , n3500 );
    and g22829 ( n1104 , n20550 , n30748 );
    not g22830 ( n7898 , n12610 );
    xor g22831 ( n2532 , n24594 , n20853 );
    xnor g22832 ( n7023 , n19089 , n20424 );
    xnor g22833 ( n8559 , n3140 , n4554 );
    or g22834 ( n4304 , n24528 , n6696 );
    and g22835 ( n10317 , n10502 , n10455 );
    not g22836 ( n18038 , n16080 );
    nor g22837 ( n31669 , n27534 , n7951 );
    and g22838 ( n14860 , n15971 , n29510 );
    nor g22839 ( n16544 , n5069 , n16108 );
    and g22840 ( n281 , n30073 , n26498 );
    and g22841 ( n17136 , n11858 , n4832 );
    not g22842 ( n16148 , n3915 );
    not g22843 ( n24192 , n23761 );
    or g22844 ( n26077 , n26657 , n7017 );
    and g22845 ( n20328 , n20099 , n18892 );
    buf g22846 ( n20865 , n1786 );
    not g22847 ( n942 , n10433 );
    and g22848 ( n27209 , n8517 , n12163 );
    xnor g22849 ( n19118 , n2251 , n14520 );
    or g22850 ( n6966 , n7158 , n10078 );
    and g22851 ( n12414 , n8128 , n14559 );
    not g22852 ( n20922 , n1195 );
    xnor g22853 ( n9697 , n12378 , n2453 );
    xnor g22854 ( n1122 , n24807 , n25699 );
    not g22855 ( n14413 , n3076 );
    not g22856 ( n5395 , n13432 );
    not g22857 ( n31425 , n19974 );
    xnor g22858 ( n25450 , n1174 , n1210 );
    nor g22859 ( n433 , n12072 , n28911 );
    xnor g22860 ( n28054 , n24184 , n15749 );
    or g22861 ( n23727 , n17255 , n5266 );
    xnor g22862 ( n18322 , n22952 , n23938 );
    not g22863 ( n9696 , n14015 );
    or g22864 ( n15339 , n28961 , n10257 );
    or g22865 ( n23328 , n16844 , n12873 );
    not g22866 ( n8524 , n22922 );
    buf g22867 ( n20427 , n23692 );
    and g22868 ( n19264 , n29540 , n6552 );
    xnor g22869 ( n24628 , n10587 , n1161 );
    or g22870 ( n21766 , n19786 , n28102 );
    not g22871 ( n4118 , n12906 );
    xnor g22872 ( n14214 , n6292 , n29831 );
    or g22873 ( n11615 , n21143 , n30235 );
    and g22874 ( n5472 , n11710 , n1632 );
    xnor g22875 ( n28065 , n30990 , n14868 );
    and g22876 ( n21683 , n18075 , n6357 );
    xnor g22877 ( n17641 , n26637 , n3715 );
    and g22878 ( n7721 , n3112 , n2133 );
    and g22879 ( n10391 , n17747 , n3974 );
    nor g22880 ( n18055 , n12711 , n2246 );
    or g22881 ( n18486 , n27247 , n2066 );
    and g22882 ( n12800 , n23264 , n29137 );
    xnor g22883 ( n12779 , n21897 , n15191 );
    not g22884 ( n5174 , n20712 );
    buf g22885 ( n28829 , n11618 );
    xnor g22886 ( n3994 , n6022 , n14171 );
    xnor g22887 ( n17284 , n25982 , n20135 );
    not g22888 ( n25637 , n19394 );
    and g22889 ( n9942 , n813 , n29090 );
    not g22890 ( n31226 , n8480 );
    xnor g22891 ( n23565 , n6502 , n23598 );
    and g22892 ( n31112 , n15932 , n2458 );
    xnor g22893 ( n30588 , n7092 , n19003 );
    or g22894 ( n24065 , n6060 , n25856 );
    or g22895 ( n24986 , n29433 , n3560 );
    xnor g22896 ( n24676 , n3537 , n21391 );
    or g22897 ( n2318 , n8988 , n4608 );
    and g22898 ( n9109 , n23733 , n22014 );
    xnor g22899 ( n3014 , n30698 , n4967 );
    xnor g22900 ( n13899 , n30777 , n21736 );
    or g22901 ( n11079 , n760 , n13878 );
    nor g22902 ( n5072 , n24510 , n11899 );
    or g22903 ( n9699 , n3297 , n9619 );
    xnor g22904 ( n18640 , n21275 , n14620 );
    or g22905 ( n10167 , n10594 , n23617 );
    and g22906 ( n18581 , n26714 , n30787 );
    not g22907 ( n23884 , n23218 );
    not g22908 ( n23554 , n28397 );
    or g22909 ( n8123 , n14035 , n6171 );
    not g22910 ( n1324 , n14473 );
    and g22911 ( n5524 , n566 , n29505 );
    not g22912 ( n990 , n6012 );
    buf g22913 ( n19701 , n18905 );
    xnor g22914 ( n10602 , n25802 , n27015 );
    nor g22915 ( n6621 , n12023 , n4340 );
    not g22916 ( n25188 , n16683 );
    xnor g22917 ( n21235 , n23046 , n16209 );
    and g22918 ( n7622 , n8069 , n24955 );
    xnor g22919 ( n21892 , n12434 , n9999 );
    not g22920 ( n18221 , n8929 );
    and g22921 ( n20698 , n1143 , n3403 );
    not g22922 ( n25995 , n31415 );
    or g22923 ( n11066 , n17852 , n21575 );
    xnor g22924 ( n5628 , n11902 , n30819 );
    or g22925 ( n2079 , n17499 , n8827 );
    and g22926 ( n4083 , n18406 , n11876 );
    or g22927 ( n8399 , n2115 , n3133 );
    xor g22928 ( n7293 , n4500 , n1025 );
    not g22929 ( n25230 , n25734 );
    or g22930 ( n505 , n15922 , n5034 );
    xnor g22931 ( n28749 , n1506 , n17133 );
    or g22932 ( n11794 , n24350 , n14785 );
    not g22933 ( n9674 , n17596 );
    xnor g22934 ( n15613 , n31485 , n19346 );
    or g22935 ( n12628 , n16986 , n28405 );
    or g22936 ( n29748 , n3894 , n9814 );
    xnor g22937 ( n9519 , n18699 , n7031 );
    xnor g22938 ( n23532 , n19092 , n11736 );
    and g22939 ( n14374 , n11242 , n35 );
    and g22940 ( n26347 , n16816 , n25526 );
    xnor g22941 ( n3340 , n14403 , n3182 );
    not g22942 ( n26377 , n24871 );
    and g22943 ( n13244 , n15576 , n21829 );
    not g22944 ( n24819 , n3138 );
    not g22945 ( n13533 , n18752 );
    xnor g22946 ( n19085 , n16809 , n22091 );
    or g22947 ( n6503 , n22619 , n24827 );
    xnor g22948 ( n4521 , n24082 , n6497 );
    not g22949 ( n17572 , n31387 );
    xnor g22950 ( n24335 , n12190 , n29287 );
    not g22951 ( n24404 , n20870 );
    xnor g22952 ( n8062 , n31354 , n3345 );
    not g22953 ( n6590 , n15971 );
    xnor g22954 ( n30821 , n6033 , n4271 );
    xnor g22955 ( n12734 , n18844 , n3956 );
    xnor g22956 ( n23254 , n28967 , n8158 );
    xnor g22957 ( n27380 , n24289 , n14690 );
    and g22958 ( n11399 , n16455 , n13610 );
    xnor g22959 ( n22140 , n23811 , n12994 );
    xnor g22960 ( n27046 , n8748 , n31146 );
    and g22961 ( n16742 , n6593 , n15295 );
    not g22962 ( n16692 , n20040 );
    and g22963 ( n30645 , n28916 , n3625 );
    not g22964 ( n17112 , n5521 );
    or g22965 ( n7089 , n1317 , n16431 );
    or g22966 ( n19560 , n31340 , n23686 );
    not g22967 ( n24865 , n9654 );
    or g22968 ( n12924 , n11859 , n24369 );
    not g22969 ( n10883 , n9500 );
    and g22970 ( n27855 , n9784 , n21099 );
    not g22971 ( n13952 , n17487 );
    nor g22972 ( n24785 , n8804 , n29084 );
    not g22973 ( n29345 , n18711 );
    and g22974 ( n26979 , n30922 , n27351 );
    or g22975 ( n9198 , n27760 , n5745 );
    xnor g22976 ( n22728 , n20950 , n23714 );
    or g22977 ( n21874 , n26583 , n7304 );
    xnor g22978 ( n25407 , n28778 , n3743 );
    and g22979 ( n16479 , n31296 , n19984 );
    and g22980 ( n29225 , n26136 , n1793 );
    or g22981 ( n19767 , n9151 , n6317 );
    or g22982 ( n3291 , n8834 , n20906 );
    xnor g22983 ( n2549 , n1466 , n9628 );
    xnor g22984 ( n492 , n10431 , n25194 );
    and g22985 ( n21886 , n11111 , n1716 );
    xnor g22986 ( n3207 , n7692 , n3106 );
    not g22987 ( n28946 , n30706 );
    not g22988 ( n23185 , n6423 );
    or g22989 ( n15287 , n29297 , n27344 );
    and g22990 ( n25223 , n14179 , n6906 );
    or g22991 ( n28405 , n9321 , n25805 );
    not g22992 ( n11810 , n23035 );
    or g22993 ( n27259 , n26203 , n7325 );
    and g22994 ( n26025 , n9383 , n21422 );
    nor g22995 ( n18705 , n28158 , n20209 );
    not g22996 ( n30161 , n27169 );
    or g22997 ( n31444 , n21542 , n4121 );
    and g22998 ( n6730 , n26757 , n8190 );
    xnor g22999 ( n18371 , n20875 , n2906 );
    or g23000 ( n10854 , n2965 , n31050 );
    nor g23001 ( n905 , n23544 , n987 );
    not g23002 ( n15256 , n24678 );
    and g23003 ( n12047 , n25087 , n14827 );
    not g23004 ( n12598 , n8838 );
    not g23005 ( n3719 , n8085 );
    not g23006 ( n20822 , n3642 );
    and g23007 ( n23974 , n14207 , n403 );
    or g23008 ( n30421 , n21597 , n14124 );
    xnor g23009 ( n12179 , n4802 , n20870 );
    xnor g23010 ( n14203 , n26532 , n2107 );
    and g23011 ( n4061 , n19082 , n13528 );
    not g23012 ( n23160 , n763 );
    xnor g23013 ( n28047 , n28607 , n11259 );
    not g23014 ( n5152 , n20307 );
    nor g23015 ( n1196 , n5638 , n11253 );
    or g23016 ( n19165 , n5631 , n14289 );
    and g23017 ( n15949 , n559 , n23770 );
    xor g23018 ( n27663 , n28498 , n28765 );
    xnor g23019 ( n14878 , n22249 , n5298 );
    or g23020 ( n7733 , n3542 , n19468 );
    not g23021 ( n4432 , n3080 );
    not g23022 ( n30464 , n5853 );
    and g23023 ( n22188 , n9055 , n8837 );
    or g23024 ( n11154 , n17089 , n20865 );
    or g23025 ( n5182 , n1819 , n11036 );
    not g23026 ( n27638 , n31366 );
    or g23027 ( n3399 , n27813 , n10361 );
    and g23028 ( n19761 , n21417 , n18071 );
    nor g23029 ( n28039 , n26255 , n14063 );
    buf g23030 ( n3677 , n24691 );
    nor g23031 ( n30204 , n3858 , n29121 );
    xnor g23032 ( n1416 , n18403 , n30405 );
    or g23033 ( n13273 , n11736 , n2628 );
    xnor g23034 ( n4736 , n18618 , n6628 );
    not g23035 ( n18113 , n10310 );
    xnor g23036 ( n24004 , n15153 , n15735 );
    xnor g23037 ( n2353 , n9043 , n9163 );
    not g23038 ( n13367 , n23131 );
    xnor g23039 ( n18112 , n4602 , n2830 );
    or g23040 ( n24859 , n2428 , n16221 );
    nor g23041 ( n25927 , n26052 , n22675 );
    or g23042 ( n21746 , n18380 , n23903 );
    not g23043 ( n9794 , n1221 );
    not g23044 ( n9569 , n12122 );
    or g23045 ( n1890 , n22514 , n24069 );
    xnor g23046 ( n30937 , n6769 , n16140 );
    xnor g23047 ( n31286 , n7237 , n17773 );
    not g23048 ( n24528 , n11611 );
    xnor g23049 ( n7797 , n3406 , n13210 );
    not g23050 ( n9523 , n4221 );
    or g23051 ( n17181 , n9411 , n19184 );
    or g23052 ( n31429 , n27064 , n4308 );
    not g23053 ( n28233 , n20365 );
    and g23054 ( n7226 , n10147 , n12315 );
    xnor g23055 ( n31763 , n9644 , n29206 );
    xnor g23056 ( n18727 , n2799 , n24464 );
    not g23057 ( n3319 , n31416 );
    and g23058 ( n14579 , n15692 , n12797 );
    and g23059 ( n25684 , n15348 , n107 );
    not g23060 ( n9327 , n15110 );
    and g23061 ( n9222 , n24693 , n26721 );
    xnor g23062 ( n22981 , n24998 , n13870 );
    not g23063 ( n1839 , n17910 );
    and g23064 ( n27998 , n25597 , n18243 );
    or g23065 ( n16589 , n23396 , n10186 );
    and g23066 ( n8539 , n5142 , n15396 );
    not g23067 ( n27065 , n18514 );
    not g23068 ( n17308 , n9653 );
    xnor g23069 ( n7386 , n31040 , n22956 );
    not g23070 ( n2882 , n12401 );
    xnor g23071 ( n28763 , n5601 , n3207 );
    and g23072 ( n13407 , n12308 , n87 );
    or g23073 ( n18847 , n6378 , n12039 );
    not g23074 ( n22151 , n8005 );
    not g23075 ( n15671 , n26771 );
    xnor g23076 ( n30256 , n21297 , n22351 );
    not g23077 ( n20178 , n315 );
    or g23078 ( n22290 , n2775 , n26763 );
    not g23079 ( n12963 , n15153 );
    not g23080 ( n8249 , n8520 );
    not g23081 ( n6121 , n2521 );
    and g23082 ( n24476 , n6221 , n30270 );
    and g23083 ( n13928 , n15404 , n12007 );
    nor g23084 ( n26527 , n1518 , n23184 );
    nor g23085 ( n4766 , n887 , n6118 );
    and g23086 ( n15953 , n7320 , n43 );
    not g23087 ( n13954 , n3383 );
    or g23088 ( n27845 , n21808 , n752 );
    or g23089 ( n8011 , n17617 , n11789 );
    or g23090 ( n28817 , n22687 , n20771 );
    not g23091 ( n7626 , n28105 );
    and g23092 ( n13937 , n10000 , n5919 );
    xnor g23093 ( n25618 , n17217 , n3182 );
    or g23094 ( n13827 , n2209 , n23166 );
    not g23095 ( n31095 , n2908 );
    xor g23096 ( n29998 , n16760 , n14356 );
    and g23097 ( n14053 , n17719 , n15566 );
    buf g23098 ( n1860 , n16563 );
    and g23099 ( n18714 , n353 , n23044 );
    and g23100 ( n29609 , n9957 , n11003 );
    not g23101 ( n9720 , n20473 );
    or g23102 ( n13778 , n10374 , n27796 );
    or g23103 ( n25501 , n29764 , n14704 );
    not g23104 ( n5876 , n24988 );
    and g23105 ( n21878 , n22511 , n4336 );
    xnor g23106 ( n26108 , n12219 , n21754 );
    and g23107 ( n14564 , n8883 , n22309 );
    or g23108 ( n22066 , n25900 , n8225 );
    not g23109 ( n10718 , n1322 );
    nor g23110 ( n27476 , n13616 , n30022 );
    xnor g23111 ( n21649 , n747 , n4632 );
    or g23112 ( n15319 , n8089 , n4683 );
    or g23113 ( n28252 , n21937 , n15599 );
    or g23114 ( n21762 , n13050 , n24340 );
    not g23115 ( n10790 , n7637 );
    and g23116 ( n24700 , n1469 , n3982 );
    not g23117 ( n23173 , n26590 );
    xnor g23118 ( n19174 , n24794 , n18955 );
    and g23119 ( n9492 , n28592 , n1552 );
    nor g23120 ( n17859 , n3668 , n11566 );
    xnor g23121 ( n4531 , n20649 , n25429 );
    or g23122 ( n30012 , n3071 , n12646 );
    xnor g23123 ( n8356 , n12884 , n16470 );
    and g23124 ( n12323 , n18856 , n6940 );
    not g23125 ( n3450 , n17270 );
    xnor g23126 ( n30856 , n19238 , n18087 );
    not g23127 ( n4014 , n26713 );
    xnor g23128 ( n19239 , n9964 , n11984 );
    or g23129 ( n30443 , n1437 , n1023 );
    xnor g23130 ( n28018 , n26902 , n29395 );
    nor g23131 ( n15880 , n4297 , n7768 );
    not g23132 ( n785 , n23960 );
    not g23133 ( n7645 , n22109 );
    xnor g23134 ( n19235 , n31443 , n22277 );
    xnor g23135 ( n25136 , n3918 , n2714 );
    xnor g23136 ( n10117 , n26789 , n19109 );
    not g23137 ( n14145 , n7187 );
    or g23138 ( n22402 , n5585 , n12141 );
    and g23139 ( n12205 , n3495 , n20023 );
    or g23140 ( n26105 , n30310 , n1440 );
    not g23141 ( n25347 , n42 );
    and g23142 ( n6000 , n3925 , n10923 );
    or g23143 ( n5048 , n4836 , n27919 );
    not g23144 ( n5032 , n2527 );
    or g23145 ( n7123 , n11294 , n14139 );
    xnor g23146 ( n21239 , n30932 , n19014 );
    or g23147 ( n1197 , n21185 , n198 );
    and g23148 ( n10294 , n28220 , n20709 );
    and g23149 ( n5837 , n14892 , n26856 );
    or g23150 ( n27328 , n655 , n13779 );
    xnor g23151 ( n5536 , n5489 , n14307 );
    nor g23152 ( n12229 , n25265 , n14446 );
    not g23153 ( n2731 , n12946 );
    not g23154 ( n362 , n24015 );
    not g23155 ( n18169 , n29028 );
    and g23156 ( n11386 , n13543 , n19017 );
    and g23157 ( n18125 , n21554 , n5224 );
    or g23158 ( n29512 , n17605 , n30338 );
    and g23159 ( n7569 , n11219 , n29344 );
    or g23160 ( n27282 , n27969 , n27652 );
    or g23161 ( n18791 , n3378 , n5504 );
    not g23162 ( n3521 , n27555 );
    not g23163 ( n8898 , n141 );
    xnor g23164 ( n25193 , n4801 , n31299 );
    or g23165 ( n5885 , n2885 , n28578 );
    xnor g23166 ( n3637 , n5472 , n13410 );
    not g23167 ( n31826 , n21647 );
    xor g23168 ( n31461 , n13985 , n30660 );
    not g23169 ( n7376 , n2978 );
    or g23170 ( n28052 , n7870 , n7263 );
    not g23171 ( n4612 , n15954 );
    or g23172 ( n4230 , n10685 , n11538 );
    not g23173 ( n28409 , n6283 );
    nor g23174 ( n21461 , n30769 , n11643 );
    or g23175 ( n9466 , n28749 , n28799 );
    nor g23176 ( n19989 , n23756 , n5246 );
    not g23177 ( n16709 , n3524 );
    or g23178 ( n31237 , n9352 , n27308 );
    xor g23179 ( n17886 , n25560 , n10064 );
    not g23180 ( n27892 , n13649 );
    xnor g23181 ( n13918 , n10426 , n29933 );
    not g23182 ( n2894 , n6449 );
    and g23183 ( n26243 , n20011 , n6980 );
    xnor g23184 ( n13150 , n24369 , n26082 );
    or g23185 ( n11221 , n12920 , n8783 );
    or g23186 ( n21745 , n23123 , n19523 );
    xnor g23187 ( n27391 , n9237 , n3396 );
    xnor g23188 ( n19094 , n6323 , n17278 );
    xnor g23189 ( n20018 , n15921 , n7115 );
    or g23190 ( n26811 , n23879 , n25846 );
    nor g23191 ( n12234 , n10291 , n20240 );
    or g23192 ( n27769 , n18585 , n28603 );
    xnor g23193 ( n15165 , n30809 , n6021 );
    not g23194 ( n28179 , n19021 );
    and g23195 ( n1341 , n11374 , n31810 );
    or g23196 ( n19267 , n18664 , n7062 );
    nor g23197 ( n27734 , n5293 , n10125 );
    and g23198 ( n18461 , n29209 , n1644 );
    and g23199 ( n13757 , n14682 , n12924 );
    not g23200 ( n11270 , n5102 );
    not g23201 ( n21568 , n10370 );
    not g23202 ( n7358 , n26683 );
    not g23203 ( n6107 , n24514 );
    nor g23204 ( n31758 , n2049 , n21711 );
    xnor g23205 ( n1276 , n6306 , n8714 );
    xnor g23206 ( n7768 , n29211 , n1613 );
    nor g23207 ( n7834 , n25518 , n26317 );
    and g23208 ( n11545 , n2582 , n16918 );
    nor g23209 ( n20683 , n15342 , n17457 );
    xnor g23210 ( n24850 , n28562 , n28983 );
    xnor g23211 ( n18882 , n24807 , n31970 );
    or g23212 ( n12417 , n20657 , n519 );
    and g23213 ( n10434 , n26843 , n25378 );
    not g23214 ( n23866 , n20643 );
    not g23215 ( n13839 , n30556 );
    xnor g23216 ( n13920 , n17582 , n14373 );
    not g23217 ( n14303 , n20791 );
    and g23218 ( n25339 , n13300 , n31060 );
    xnor g23219 ( n20358 , n28781 , n18165 );
    and g23220 ( n26895 , n22879 , n28123 );
    xnor g23221 ( n11815 , n16820 , n4448 );
    and g23222 ( n12458 , n6518 , n28664 );
    buf g23223 ( n11740 , n28135 );
    or g23224 ( n20840 , n2046 , n8814 );
    xnor g23225 ( n7799 , n25607 , n10626 );
    not g23226 ( n15201 , n12018 );
    xnor g23227 ( n30263 , n28538 , n21728 );
    not g23228 ( n9941 , n9266 );
    not g23229 ( n29497 , n13674 );
    xnor g23230 ( n12587 , n8761 , n17287 );
    nor g23231 ( n20810 , n29063 , n19268 );
    xnor g23232 ( n31721 , n4688 , n16561 );
    and g23233 ( n23680 , n19028 , n30589 );
    or g23234 ( n13823 , n22867 , n12030 );
    and g23235 ( n14198 , n13081 , n23342 );
    not g23236 ( n31191 , n10602 );
    nor g23237 ( n11189 , n30326 , n29153 );
    not g23238 ( n19678 , n5572 );
    and g23239 ( n8765 , n29935 , n16952 );
    nor g23240 ( n26912 , n5614 , n29791 );
    not g23241 ( n30040 , n7588 );
    and g23242 ( n4534 , n30549 , n6874 );
    not g23243 ( n23651 , n11679 );
    nor g23244 ( n8025 , n10893 , n22447 );
    or g23245 ( n4373 , n17240 , n3273 );
    xnor g23246 ( n15715 , n27535 , n5559 );
    or g23247 ( n25309 , n4273 , n15199 );
    or g23248 ( n2142 , n24573 , n5511 );
    or g23249 ( n23961 , n30245 , n22005 );
    not g23250 ( n9108 , n17866 );
    or g23251 ( n18171 , n14 , n26550 );
    xnor g23252 ( n25911 , n31070 , n29293 );
    or g23253 ( n26613 , n27072 , n4 );
    not g23254 ( n31498 , n21375 );
    and g23255 ( n30693 , n15907 , n16173 );
    and g23256 ( n3193 , n31961 , n1312 );
    or g23257 ( n10659 , n28697 , n20313 );
    not g23258 ( n903 , n24425 );
    xnor g23259 ( n13970 , n13998 , n28397 );
    or g23260 ( n9755 , n18963 , n24996 );
    xnor g23261 ( n28892 , n23359 , n11110 );
    xnor g23262 ( n19396 , n29543 , n6356 );
    xnor g23263 ( n30741 , n28876 , n2055 );
    and g23264 ( n16657 , n30176 , n22104 );
    xnor g23265 ( n1515 , n9827 , n1358 );
    and g23266 ( n25520 , n25353 , n25343 );
    not g23267 ( n14920 , n3884 );
    not g23268 ( n22129 , n18529 );
    or g23269 ( n4461 , n16017 , n17288 );
    not g23270 ( n7638 , n1867 );
    and g23271 ( n31031 , n9819 , n18626 );
    xnor g23272 ( n5916 , n14882 , n24008 );
    xnor g23273 ( n6280 , n29383 , n2810 );
    not g23274 ( n30303 , n15586 );
    nor g23275 ( n30646 , n5559 , n6836 );
    and g23276 ( n9028 , n21678 , n22280 );
    or g23277 ( n918 , n11171 , n20999 );
    and g23278 ( n30304 , n15837 , n13183 );
    not g23279 ( n3438 , n11064 );
    not g23280 ( n20030 , n8369 );
    and g23281 ( n13821 , n30428 , n1417 );
    not g23282 ( n2282 , n51 );
    not g23283 ( n9220 , n15335 );
    not g23284 ( n8612 , n5781 );
    or g23285 ( n22941 , n20347 , n29218 );
    not g23286 ( n28438 , n16655 );
    xnor g23287 ( n26906 , n29153 , n2610 );
    xor g23288 ( n9099 , n20991 , n6558 );
    xnor g23289 ( n31575 , n19163 , n12327 );
    xnor g23290 ( n10168 , n13632 , n19791 );
    not g23291 ( n11143 , n7011 );
    or g23292 ( n21403 , n16161 , n29674 );
    xnor g23293 ( n25666 , n7414 , n3080 );
    or g23294 ( n8190 , n31889 , n5697 );
    or g23295 ( n18064 , n10595 , n7440 );
    xnor g23296 ( n21469 , n18056 , n24800 );
    not g23297 ( n18258 , n7083 );
    xnor g23298 ( n9418 , n8883 , n23758 );
    xnor g23299 ( n18266 , n10486 , n19811 );
    not g23300 ( n20804 , n1532 );
    and g23301 ( n26862 , n13717 , n27595 );
    and g23302 ( n14253 , n7733 , n13246 );
    xnor g23303 ( n12728 , n15661 , n28587 );
    not g23304 ( n11236 , n12566 );
    not g23305 ( n5407 , n7433 );
    nor g23306 ( n2756 , n256 , n29950 );
    or g23307 ( n11275 , n20632 , n30530 );
    not g23308 ( n11543 , n3475 );
    and g23309 ( n3143 , n5539 , n3152 );
    xnor g23310 ( n1447 , n26582 , n3590 );
    xnor g23311 ( n1592 , n1193 , n11482 );
    not g23312 ( n9467 , n31942 );
    not g23313 ( n6839 , n9935 );
    not g23314 ( n5542 , n7078 );
    or g23315 ( n10935 , n17585 , n3101 );
    not g23316 ( n12397 , n23339 );
    or g23317 ( n18732 , n6472 , n3519 );
    and g23318 ( n22682 , n24810 , n13051 );
    not g23319 ( n23634 , n31366 );
    or g23320 ( n3003 , n26598 , n31806 );
    xnor g23321 ( n28161 , n3259 , n2883 );
    and g23322 ( n30376 , n28495 , n22790 );
    or g23323 ( n5344 , n13454 , n30458 );
    and g23324 ( n21944 , n15103 , n19860 );
    xnor g23325 ( n16081 , n26076 , n5247 );
    xnor g23326 ( n11354 , n5097 , n29365 );
    or g23327 ( n25313 , n13162 , n12857 );
    not g23328 ( n12640 , n3058 );
    or g23329 ( n13898 , n29226 , n4079 );
    or g23330 ( n20948 , n19054 , n12441 );
    and g23331 ( n5302 , n20886 , n24984 );
    or g23332 ( n15442 , n19890 , n7769 );
    not g23333 ( n14693 , n25566 );
    or g23334 ( n7510 , n15467 , n23408 );
    and g23335 ( n737 , n18834 , n31946 );
    nor g23336 ( n6568 , n29145 , n12955 );
    xnor g23337 ( n1933 , n2977 , n13540 );
    not g23338 ( n23750 , n5202 );
    not g23339 ( n16865 , n7010 );
    not g23340 ( n31705 , n2461 );
    not g23341 ( n14370 , n26198 );
    or g23342 ( n22817 , n26699 , n27685 );
    not g23343 ( n61 , n12953 );
    or g23344 ( n8719 , n6888 , n30617 );
    not g23345 ( n4154 , n731 );
    or g23346 ( n15688 , n24917 , n25689 );
    or g23347 ( n3431 , n27147 , n15510 );
    or g23348 ( n1013 , n10628 , n30397 );
    not g23349 ( n16688 , n15335 );
    or g23350 ( n28842 , n18202 , n11466 );
    xnor g23351 ( n25306 , n18273 , n2964 );
    not g23352 ( n24552 , n22710 );
    and g23353 ( n25287 , n21178 , n283 );
    and g23354 ( n13896 , n23830 , n29232 );
    xnor g23355 ( n27849 , n11017 , n25012 );
    xnor g23356 ( n17530 , n26129 , n25549 );
    or g23357 ( n17800 , n9655 , n2794 );
    and g23358 ( n25955 , n22648 , n22992 );
    or g23359 ( n16165 , n17867 , n26905 );
    xnor g23360 ( n23732 , n18850 , n23047 );
    xnor g23361 ( n18731 , n10762 , n2460 );
    or g23362 ( n8429 , n29200 , n18069 );
    not g23363 ( n719 , n24118 );
    and g23364 ( n26482 , n17785 , n20681 );
    not g23365 ( n19643 , n6249 );
    not g23366 ( n28940 , n9367 );
    nor g23367 ( n872 , n4350 , n22371 );
    or g23368 ( n103 , n18754 , n31328 );
    and g23369 ( n3180 , n18732 , n2758 );
    not g23370 ( n7420 , n6240 );
    not g23371 ( n20467 , n2054 );
    and g23372 ( n8830 , n28406 , n18187 );
    not g23373 ( n16836 , n21252 );
    xnor g23374 ( n11994 , n3643 , n154 );
    xnor g23375 ( n25295 , n23224 , n17720 );
    or g23376 ( n20645 , n17331 , n27723 );
    not g23377 ( n24414 , n8698 );
    not g23378 ( n10859 , n8516 );
    not g23379 ( n3213 , n13710 );
    and g23380 ( n16179 , n207 , n28743 );
    not g23381 ( n19649 , n16301 );
    nor g23382 ( n26551 , n1692 , n11643 );
    not g23383 ( n11587 , n13065 );
    or g23384 ( n23325 , n17699 , n1223 );
    xnor g23385 ( n6258 , n18841 , n10674 );
    not g23386 ( n12739 , n9135 );
    and g23387 ( n4029 , n3111 , n27050 );
    and g23388 ( n29937 , n19644 , n21222 );
    not g23389 ( n10379 , n22723 );
    or g23390 ( n1185 , n29877 , n6806 );
    or g23391 ( n28214 , n6803 , n2736 );
    xnor g23392 ( n26932 , n8665 , n9805 );
    buf g23393 ( n24129 , n6056 );
    xnor g23394 ( n31695 , n29504 , n6274 );
    xnor g23395 ( n12031 , n19804 , n10914 );
    or g23396 ( n12875 , n29022 , n18659 );
    or g23397 ( n16341 , n141 , n27853 );
    or g23398 ( n18290 , n6354 , n18609 );
    xnor g23399 ( n864 , n7498 , n28671 );
    xnor g23400 ( n14655 , n8871 , n26877 );
    or g23401 ( n6723 , n29822 , n4552 );
    not g23402 ( n27461 , n5037 );
    and g23403 ( n20930 , n20496 , n16458 );
    not g23404 ( n1473 , n826 );
    or g23405 ( n13691 , n11478 , n11648 );
    xnor g23406 ( n26604 , n25856 , n21597 );
    xnor g23407 ( n9608 , n2158 , n7511 );
    or g23408 ( n28529 , n21104 , n22907 );
    not g23409 ( n880 , n12566 );
    not g23410 ( n10891 , n31250 );
    or g23411 ( n13861 , n28947 , n12742 );
    xnor g23412 ( n28918 , n6549 , n12030 );
    and g23413 ( n29893 , n15461 , n6771 );
    or g23414 ( n20847 , n17983 , n257 );
    or g23415 ( n7618 , n5480 , n1668 );
    or g23416 ( n1486 , n26449 , n12829 );
    not g23417 ( n30384 , n11322 );
    nor g23418 ( n2766 , n19125 , n12664 );
    or g23419 ( n5138 , n21660 , n1490 );
    not g23420 ( n20728 , n2483 );
    xnor g23421 ( n3678 , n12258 , n5805 );
    not g23422 ( n11416 , n9820 );
    and g23423 ( n13541 , n13881 , n20036 );
    not g23424 ( n26438 , n13859 );
    xnor g23425 ( n29208 , n27200 , n5133 );
    or g23426 ( n13731 , n19720 , n18345 );
    nor g23427 ( n30230 , n2231 , n9720 );
    xor g23428 ( n30360 , n26217 , n22866 );
    xnor g23429 ( n17497 , n16325 , n6192 );
    nor g23430 ( n3075 , n10050 , n15398 );
    or g23431 ( n1399 , n14324 , n3461 );
    and g23432 ( n22975 , n26946 , n4962 );
    nor g23433 ( n14765 , n24681 , n15341 );
    or g23434 ( n28190 , n11046 , n31588 );
    and g23435 ( n17446 , n7844 , n29444 );
    and g23436 ( n24685 , n7073 , n4395 );
    not g23437 ( n28987 , n9645 );
    and g23438 ( n10857 , n5078 , n14992 );
    xnor g23439 ( n16450 , n30433 , n12221 );
    and g23440 ( n16354 , n7622 , n5691 );
    and g23441 ( n21840 , n9385 , n14216 );
    or g23442 ( n31605 , n14914 , n26357 );
    not g23443 ( n13321 , n4188 );
    xnor g23444 ( n1481 , n6947 , n8336 );
    or g23445 ( n21460 , n6093 , n14223 );
    not g23446 ( n1889 , n15320 );
    xnor g23447 ( n15257 , n25082 , n10693 );
    buf g23448 ( n24784 , n7044 );
    not g23449 ( n11820 , n29854 );
    or g23450 ( n25975 , n13476 , n14724 );
    not g23451 ( n11630 , n11889 );
    not g23452 ( n7901 , n28021 );
    or g23453 ( n7653 , n9024 , n22768 );
    xnor g23454 ( n23799 , n9 , n30688 );
    or g23455 ( n4321 , n13549 , n30703 );
    not g23456 ( n2971 , n3602 );
    or g23457 ( n10896 , n5071 , n5924 );
    not g23458 ( n31960 , n26353 );
    xnor g23459 ( n24223 , n15408 , n15936 );
    not g23460 ( n24130 , n31960 );
    xnor g23461 ( n3190 , n29238 , n1095 );
    and g23462 ( n23608 , n12826 , n30466 );
    or g23463 ( n24370 , n11014 , n24125 );
    xor g23464 ( n29361 , n14274 , n4836 );
    or g23465 ( n8169 , n10523 , n339 );
    not g23466 ( n1807 , n19704 );
    and g23467 ( n3894 , n12841 , n23023 );
    xnor g23468 ( n27660 , n31359 , n12679 );
    or g23469 ( n6119 , n1942 , n5483 );
    or g23470 ( n3768 , n10955 , n3701 );
    xnor g23471 ( n27587 , n28310 , n1066 );
    not g23472 ( n25324 , n858 );
    not g23473 ( n20842 , n5358 );
    not g23474 ( n25458 , n9480 );
    xnor g23475 ( n12737 , n2647 , n26524 );
    and g23476 ( n19111 , n5855 , n17520 );
    xnor g23477 ( n12561 , n3181 , n1960 );
    xnor g23478 ( n12153 , n1855 , n30829 );
    and g23479 ( n25167 , n20056 , n21272 );
    xnor g23480 ( n25058 , n8991 , n31204 );
    or g23481 ( n1323 , n31403 , n7199 );
    and g23482 ( n13650 , n3834 , n30796 );
    xnor g23483 ( n618 , n20458 , n18985 );
    not g23484 ( n16772 , n14269 );
    and g23485 ( n30610 , n20203 , n21654 );
    xnor g23486 ( n28609 , n7301 , n3951 );
    not g23487 ( n27441 , n12251 );
    xnor g23488 ( n5400 , n27811 , n20238 );
    xnor g23489 ( n21981 , n5729 , n12253 );
    or g23490 ( n12655 , n8497 , n31805 );
    xnor g23491 ( n14699 , n24215 , n23170 );
    not g23492 ( n18744 , n28999 );
    xnor g23493 ( n5212 , n7693 , n26542 );
    not g23494 ( n23879 , n21291 );
    xnor g23495 ( n8051 , n22742 , n3599 );
    not g23496 ( n17123 , n13693 );
    xnor g23497 ( n2381 , n26825 , n19720 );
    or g23498 ( n20003 , n24467 , n7321 );
    or g23499 ( n23399 , n19629 , n21625 );
    or g23500 ( n13070 , n11897 , n22333 );
    or g23501 ( n10273 , n27793 , n30851 );
    and g23502 ( n30488 , n25609 , n21511 );
    not g23503 ( n13599 , n16291 );
    xnor g23504 ( n19183 , n5263 , n26860 );
    xnor g23505 ( n1161 , n10980 , n20525 );
    nor g23506 ( n11105 , n22203 , n5181 );
    buf g23507 ( n4451 , n5576 );
    xnor g23508 ( n8043 , n652 , n23775 );
    xnor g23509 ( n7435 , n14637 , n21262 );
    xnor g23510 ( n14259 , n22061 , n8090 );
    or g23511 ( n12855 , n25115 , n7229 );
    and g23512 ( n31794 , n2946 , n11809 );
    or g23513 ( n28255 , n4005 , n4637 );
    xnor g23514 ( n13570 , n29368 , n25242 );
    xnor g23515 ( n22180 , n31436 , n30865 );
    not g23516 ( n5940 , n10862 );
    not g23517 ( n17294 , n8509 );
    or g23518 ( n10590 , n926 , n16936 );
    or g23519 ( n28519 , n6326 , n13951 );
    or g23520 ( n9516 , n8860 , n19834 );
    not g23521 ( n21487 , n6300 );
    and g23522 ( n12884 , n24292 , n28848 );
    not g23523 ( n25026 , n3514 );
    and g23524 ( n12137 , n17453 , n22465 );
    not g23525 ( n30733 , n4287 );
    xnor g23526 ( n22408 , n11408 , n10506 );
    xnor g23527 ( n25208 , n6308 , n28661 );
    not g23528 ( n1238 , n21508 );
    and g23529 ( n15972 , n21812 , n9348 );
    xnor g23530 ( n4276 , n28315 , n26598 );
    xnor g23531 ( n14822 , n7877 , n29565 );
    not g23532 ( n29168 , n22216 );
    not g23533 ( n22094 , n28170 );
    nor g23534 ( n19485 , n23960 , n12293 );
    nor g23535 ( n13213 , n25579 , n25189 );
    or g23536 ( n24354 , n23368 , n4950 );
    not g23537 ( n25383 , n16987 );
    xnor g23538 ( n11708 , n24923 , n16007 );
    not g23539 ( n10133 , n19632 );
    not g23540 ( n13020 , n15906 );
    not g23541 ( n13579 , n1692 );
    and g23542 ( n17700 , n20960 , n9316 );
    and g23543 ( n5286 , n8588 , n10808 );
    and g23544 ( n28379 , n19197 , n22090 );
    not g23545 ( n21435 , n27716 );
    and g23546 ( n31936 , n2151 , n19164 );
    not g23547 ( n8440 , n6840 );
    not g23548 ( n2294 , n5187 );
    and g23549 ( n5155 , n17654 , n22433 );
    and g23550 ( n19899 , n27707 , n7038 );
    xnor g23551 ( n9891 , n29098 , n17853 );
    and g23552 ( n27428 , n16046 , n4596 );
    not g23553 ( n18585 , n13414 );
    and g23554 ( n19351 , n4385 , n3965 );
    xnor g23555 ( n3730 , n11658 , n19132 );
    not g23556 ( n17454 , n29493 );
    xnor g23557 ( n21563 , n31236 , n30588 );
    or g23558 ( n18521 , n21286 , n30105 );
    or g23559 ( n11013 , n10334 , n7046 );
    xnor g23560 ( n1283 , n1334 , n12951 );
    xor g23561 ( n3063 , n19533 , n5012 );
    and g23562 ( n2181 , n22173 , n16851 );
    and g23563 ( n16721 , n777 , n8005 );
    not g23564 ( n6391 , n914 );
    or g23565 ( n19576 , n18002 , n24280 );
    not g23566 ( n20176 , n11071 );
    or g23567 ( n23073 , n3193 , n2874 );
    not g23568 ( n5791 , n12301 );
    not g23569 ( n6216 , n5573 );
    or g23570 ( n4017 , n12330 , n19201 );
    or g23571 ( n31542 , n28786 , n23263 );
    not g23572 ( n15341 , n12375 );
    and g23573 ( n2297 , n28076 , n11768 );
    not g23574 ( n351 , n23523 );
    not g23575 ( n6867 , n10404 );
    and g23576 ( n25250 , n29973 , n29465 );
    xnor g23577 ( n22656 , n31205 , n30326 );
    or g23578 ( n17980 , n9604 , n24522 );
    xnor g23579 ( n26037 , n10289 , n6399 );
    not g23580 ( n22363 , n25208 );
    not g23581 ( n19864 , n6620 );
    nor g23582 ( n5223 , n6005 , n7858 );
    or g23583 ( n29350 , n960 , n10396 );
    xnor g23584 ( n16007 , n19010 , n10643 );
    not g23585 ( n15934 , n2462 );
    xnor g23586 ( n26051 , n26655 , n17255 );
    not g23587 ( n26533 , n10742 );
    or g23588 ( n3088 , n12828 , n2977 );
    and g23589 ( n28955 , n953 , n5240 );
    xnor g23590 ( n25432 , n20140 , n14964 );
    xor g23591 ( n3873 , n3762 , n14419 );
    and g23592 ( n5403 , n2841 , n28667 );
    not g23593 ( n26825 , n30997 );
    xnor g23594 ( n5008 , n18091 , n7882 );
    not g23595 ( n29010 , n30089 );
    xnor g23596 ( n4149 , n27567 , n8427 );
    not g23597 ( n31467 , n22184 );
    xnor g23598 ( n17749 , n20155 , n14624 );
    or g23599 ( n19644 , n2926 , n19944 );
    xor g23600 ( n12178 , n6573 , n18528 );
    not g23601 ( n8092 , n22184 );
    xnor g23602 ( n11388 , n4612 , n9638 );
    xnor g23603 ( n16888 , n31025 , n21981 );
    xor g23604 ( n28531 , n23722 , n31900 );
    not g23605 ( n28260 , n13604 );
    not g23606 ( n20567 , n13044 );
    xnor g23607 ( n18161 , n12294 , n31863 );
    or g23608 ( n4651 , n12658 , n17727 );
    or g23609 ( n30437 , n22745 , n16839 );
    or g23610 ( n14594 , n667 , n25735 );
    not g23611 ( n23197 , n30074 );
    and g23612 ( n21578 , n24780 , n22740 );
    and g23613 ( n12969 , n3445 , n16841 );
    xnor g23614 ( n19233 , n13 , n5736 );
    not g23615 ( n25536 , n11498 );
    and g23616 ( n27024 , n30450 , n19588 );
    not g23617 ( n25320 , n4374 );
    xnor g23618 ( n28891 , n2218 , n25291 );
    and g23619 ( n11046 , n13155 , n28642 );
    not g23620 ( n20569 , n20428 );
    xnor g23621 ( n3019 , n13924 , n14938 );
    not g23622 ( n24926 , n27696 );
    not g23623 ( n3904 , n17798 );
    or g23624 ( n2306 , n9740 , n6149 );
    or g23625 ( n25216 , n28845 , n8436 );
    nor g23626 ( n2624 , n29249 , n30546 );
    xor g23627 ( n7174 , n13279 , n14228 );
    xnor g23628 ( n2595 , n913 , n26791 );
    nor g23629 ( n7577 , n23124 , n22282 );
    and g23630 ( n11089 , n14165 , n16176 );
    nor g23631 ( n31521 , n2139 , n3085 );
    not g23632 ( n28177 , n12242 );
    and g23633 ( n19763 , n8391 , n7447 );
    nor g23634 ( n8668 , n25809 , n6826 );
    xnor g23635 ( n30085 , n19209 , n1676 );
    or g23636 ( n2265 , n15708 , n7026 );
    not g23637 ( n18098 , n16214 );
    not g23638 ( n2778 , n7988 );
    not g23639 ( n2469 , n4330 );
    not g23640 ( n7669 , n3620 );
    nor g23641 ( n3451 , n17368 , n26686 );
    and g23642 ( n27914 , n10366 , n9064 );
    or g23643 ( n28209 , n11540 , n20787 );
    xor g23644 ( n1677 , n11824 , n26846 );
    or g23645 ( n28439 , n24139 , n11879 );
    nor g23646 ( n3670 , n7241 , n17798 );
    and g23647 ( n29044 , n9932 , n27208 );
    or g23648 ( n7599 , n14900 , n30316 );
    or g23649 ( n558 , n28241 , n24369 );
    or g23650 ( n15868 , n9567 , n11280 );
    or g23651 ( n11768 , n29727 , n23819 );
    and g23652 ( n6167 , n31599 , n1486 );
    or g23653 ( n8833 , n5205 , n28447 );
    xnor g23654 ( n2167 , n19655 , n2405 );
    xnor g23655 ( n24899 , n5111 , n18612 );
    xnor g23656 ( n24224 , n21104 , n2798 );
    xnor g23657 ( n29938 , n21619 , n20455 );
    and g23658 ( n20378 , n3334 , n3291 );
    not g23659 ( n17176 , n26072 );
    nor g23660 ( n9306 , n1696 , n24149 );
    or g23661 ( n21596 , n1051 , n26482 );
    or g23662 ( n13408 , n23955 , n31861 );
    and g23663 ( n24054 , n12571 , n26976 );
    nor g23664 ( n27779 , n30998 , n10120 );
    or g23665 ( n22735 , n17355 , n8477 );
    or g23666 ( n21296 , n1759 , n4909 );
    not g23667 ( n4312 , n192 );
    or g23668 ( n2902 , n10021 , n8277 );
    xnor g23669 ( n27344 , n11044 , n10231 );
    and g23670 ( n10281 , n18600 , n14240 );
    nor g23671 ( n20744 , n21184 , n19836 );
    or g23672 ( n26434 , n24413 , n10230 );
    and g23673 ( n7617 , n4068 , n17666 );
    or g23674 ( n25379 , n22665 , n20815 );
    not g23675 ( n18491 , n19512 );
    not g23676 ( n21824 , n3765 );
    nor g23677 ( n22608 , n9414 , n20906 );
    and g23678 ( n4756 , n27821 , n9197 );
    not g23679 ( n27908 , n23767 );
    or g23680 ( n17865 , n14704 , n19820 );
    or g23681 ( n9083 , n22434 , n30691 );
    not g23682 ( n5765 , n27441 );
    not g23683 ( n15448 , n23508 );
    or g23684 ( n8128 , n15560 , n24813 );
    xnor g23685 ( n16951 , n29760 , n10797 );
    not g23686 ( n11181 , n3535 );
    or g23687 ( n30920 , n30532 , n13214 );
    nor g23688 ( n24178 , n18063 , n4834 );
    and g23689 ( n20498 , n19645 , n11758 );
    and g23690 ( n30970 , n8052 , n10835 );
    not g23691 ( n17261 , n26948 );
    or g23692 ( n27990 , n29938 , n3332 );
    nor g23693 ( n1825 , n10450 , n16144 );
    or g23694 ( n722 , n1329 , n6571 );
    xnor g23695 ( n21260 , n24161 , n15492 );
    nor g23696 ( n6788 , n26763 , n27175 );
    or g23697 ( n13721 , n12504 , n19729 );
    or g23698 ( n18152 , n22609 , n12387 );
    or g23699 ( n3760 , n25644 , n29534 );
    or g23700 ( n30764 , n7476 , n6781 );
    not g23701 ( n21660 , n23122 );
    xnor g23702 ( n11576 , n2683 , n22416 );
    and g23703 ( n123 , n3191 , n27126 );
    xnor g23704 ( n24649 , n12215 , n23992 );
    or g23705 ( n3813 , n9544 , n19806 );
    and g23706 ( n7331 , n10561 , n26661 );
    or g23707 ( n15434 , n17570 , n16129 );
    not g23708 ( n6578 , n666 );
    and g23709 ( n18689 , n20618 , n27369 );
    or g23710 ( n4989 , n11524 , n31959 );
    not g23711 ( n4133 , n8826 );
    nor g23712 ( n21872 , n23996 , n4868 );
    not g23713 ( n20748 , n16113 );
    and g23714 ( n15626 , n28130 , n25052 );
    or g23715 ( n18141 , n9033 , n27379 );
    or g23716 ( n2972 , n1830 , n31638 );
    not g23717 ( n28499 , n9373 );
    not g23718 ( n10931 , n19492 );
    or g23719 ( n5589 , n31192 , n16766 );
    or g23720 ( n9231 , n8310 , n7249 );
    not g23721 ( n995 , n1260 );
    not g23722 ( n2178 , n19466 );
    xnor g23723 ( n5782 , n16570 , n16785 );
    xnor g23724 ( n20159 , n8800 , n6882 );
    or g23725 ( n1081 , n8295 , n30298 );
    or g23726 ( n31594 , n21180 , n8816 );
    xnor g23727 ( n7190 , n22497 , n12971 );
    or g23728 ( n19045 , n10354 , n649 );
    not g23729 ( n1037 , n5935 );
    not g23730 ( n23738 , n23503 );
    not g23731 ( n8662 , n30720 );
    and g23732 ( n13592 , n26126 , n2838 );
    and g23733 ( n23616 , n26463 , n22473 );
    and g23734 ( n17292 , n1215 , n11099 );
    and g23735 ( n26367 , n17675 , n11248 );
    and g23736 ( n10697 , n2223 , n30960 );
    and g23737 ( n5871 , n8350 , n2495 );
    and g23738 ( n28240 , n9060 , n15392 );
    xnor g23739 ( n26269 , n21578 , n20767 );
    xnor g23740 ( n22164 , n8032 , n23516 );
    xnor g23741 ( n28141 , n31909 , n3999 );
    or g23742 ( n22662 , n21644 , n31402 );
    xnor g23743 ( n18792 , n9112 , n8456 );
    or g23744 ( n26035 , n10602 , n4344 );
    not g23745 ( n21273 , n2358 );
    or g23746 ( n22249 , n3242 , n15093 );
    and g23747 ( n22768 , n4411 , n11224 );
    not g23748 ( n2741 , n22591 );
    not g23749 ( n8739 , n20832 );
    nor g23750 ( n17727 , n1609 , n12800 );
    not g23751 ( n31500 , n30831 );
    nor g23752 ( n25635 , n3863 , n1238 );
    nor g23753 ( n11441 , n3548 , n14735 );
    nor g23754 ( n11304 , n29615 , n1488 );
    xnor g23755 ( n29790 , n20715 , n28638 );
    and g23756 ( n17614 , n19719 , n19947 );
    not g23757 ( n27470 , n21466 );
    nor g23758 ( n28676 , n24068 , n15081 );
    not g23759 ( n28490 , n16059 );
    not g23760 ( n29867 , n32032 );
    xnor g23761 ( n24383 , n28665 , n14576 );
    xnor g23762 ( n9400 , n31725 , n17910 );
    xnor g23763 ( n7363 , n27745 , n17947 );
    xnor g23764 ( n4297 , n17232 , n24005 );
    xnor g23765 ( n1096 , n14558 , n25760 );
    not g23766 ( n10785 , n8326 );
    xnor g23767 ( n9497 , n6094 , n23378 );
    or g23768 ( n1664 , n624 , n19298 );
    not g23769 ( n12475 , n26658 );
    and g23770 ( n29230 , n28889 , n686 );
    and g23771 ( n22612 , n18956 , n8062 );
    and g23772 ( n5318 , n10160 , n15879 );
    xnor g23773 ( n16652 , n13513 , n25057 );
    or g23774 ( n20193 , n14711 , n19803 );
    xnor g23775 ( n8575 , n8288 , n12063 );
    or g23776 ( n20814 , n22143 , n26951 );
    xnor g23777 ( n297 , n30264 , n15877 );
    not g23778 ( n29320 , n16269 );
    or g23779 ( n15590 , n29751 , n4238 );
    or g23780 ( n1373 , n22855 , n12788 );
    xnor g23781 ( n28765 , n21102 , n16609 );
    nor g23782 ( n25282 , n31676 , n12195 );
    not g23783 ( n12459 , n22020 );
    and g23784 ( n28037 , n1330 , n15084 );
    xnor g23785 ( n31837 , n9396 , n9948 );
    xnor g23786 ( n29494 , n6402 , n9588 );
    not g23787 ( n16784 , n18136 );
    or g23788 ( n10495 , n19738 , n13003 );
    and g23789 ( n22671 , n17919 , n22163 );
    or g23790 ( n28759 , n2514 , n13592 );
    nor g23791 ( n21077 , n5963 , n5561 );
    and g23792 ( n13820 , n9853 , n6267 );
    not g23793 ( n27345 , n16732 );
    or g23794 ( n22128 , n8988 , n23094 );
    or g23795 ( n17758 , n12207 , n12931 );
    or g23796 ( n12419 , n2665 , n7548 );
    not g23797 ( n31718 , n1923 );
    xnor g23798 ( n725 , n27504 , n4844 );
    or g23799 ( n20688 , n19460 , n17636 );
    or g23800 ( n21251 , n22045 , n23202 );
    or g23801 ( n7366 , n12764 , n2071 );
    or g23802 ( n31776 , n3028 , n24856 );
    and g23803 ( n20879 , n7691 , n12289 );
    not g23804 ( n29384 , n8289 );
    or g23805 ( n25184 , n30943 , n31710 );
    xnor g23806 ( n25860 , n11623 , n29303 );
    xnor g23807 ( n15790 , n19560 , n9774 );
    or g23808 ( n12517 , n4595 , n12264 );
    and g23809 ( n17988 , n30192 , n2647 );
    and g23810 ( n15120 , n29742 , n3777 );
    xnor g23811 ( n22794 , n15298 , n19534 );
    or g23812 ( n29334 , n12062 , n9907 );
    or g23813 ( n18740 , n2953 , n7912 );
    xnor g23814 ( n1424 , n4338 , n5228 );
    not g23815 ( n4211 , n20026 );
    xor g23816 ( n19857 , n28851 , n25796 );
    or g23817 ( n30325 , n31490 , n2362 );
    xnor g23818 ( n6313 , n27855 , n30390 );
    nor g23819 ( n3577 , n27761 , n21833 );
    xnor g23820 ( n21998 , n22890 , n12807 );
    xor g23821 ( n9502 , n22139 , n18203 );
    and g23822 ( n8351 , n22078 , n28908 );
    buf g23823 ( n16061 , n804 );
    not g23824 ( n20158 , n23813 );
    and g23825 ( n19714 , n22520 , n24189 );
    xnor g23826 ( n118 , n22926 , n19841 );
    not g23827 ( n197 , n18657 );
    xnor g23828 ( n20385 , n19519 , n9182 );
    nor g23829 ( n17274 , n25687 , n11178 );
    or g23830 ( n15047 , n27534 , n13725 );
    nor g23831 ( n8340 , n24137 , n10133 );
    not g23832 ( n27910 , n23100 );
    nor g23833 ( n7613 , n3490 , n23597 );
    nor g23834 ( n17689 , n12987 , n16843 );
    or g23835 ( n27794 , n14538 , n21855 );
    xor g23836 ( n5562 , n10525 , n6888 );
    nor g23837 ( n16212 , n7379 , n16076 );
    not g23838 ( n22238 , n5531 );
    not g23839 ( n31032 , n6276 );
    not g23840 ( n8848 , n7160 );
    xnor g23841 ( n9168 , n21988 , n20418 );
    not g23842 ( n19705 , n9061 );
    or g23843 ( n15477 , n17736 , n24054 );
    not g23844 ( n22736 , n16998 );
    not g23845 ( n30632 , n7593 );
    not g23846 ( n1415 , n18098 );
    and g23847 ( n28769 , n7831 , n4304 );
    or g23848 ( n28536 , n15008 , n22006 );
    nor g23849 ( n2658 , n20067 , n9824 );
    or g23850 ( n480 , n5594 , n7488 );
    or g23851 ( n24112 , n28503 , n29354 );
    nor g23852 ( n8310 , n963 , n26362 );
    xnor g23853 ( n1967 , n10922 , n21249 );
    or g23854 ( n29953 , n13838 , n25152 );
    or g23855 ( n22556 , n26034 , n11904 );
    or g23856 ( n5978 , n19255 , n23676 );
    or g23857 ( n16423 , n14981 , n16303 );
    not g23858 ( n22528 , n22512 );
    nor g23859 ( n16407 , n3863 , n18184 );
    or g23860 ( n25799 , n29427 , n21130 );
    or g23861 ( n24410 , n20683 , n13633 );
    not g23862 ( n7891 , n4347 );
    and g23863 ( n21935 , n5100 , n19756 );
    and g23864 ( n29438 , n9261 , n10809 );
    or g23865 ( n19990 , n21871 , n4033 );
    xor g23866 ( n21561 , n11923 , n12322 );
    or g23867 ( n1085 , n25195 , n18034 );
    xnor g23868 ( n5029 , n15386 , n17691 );
    not g23869 ( n27163 , n25001 );
    or g23870 ( n31154 , n26716 , n5913 );
    not g23871 ( n7256 , n1685 );
    not g23872 ( n25376 , n12926 );
    and g23873 ( n7679 , n21126 , n30421 );
    nor g23874 ( n19313 , n29466 , n16688 );
    and g23875 ( n9199 , n20244 , n24233 );
    not g23876 ( n6273 , n17517 );
    and g23877 ( n8831 , n31923 , n22835 );
    xnor g23878 ( n7809 , n21963 , n23934 );
    not g23879 ( n8846 , n11880 );
    and g23880 ( n13024 , n786 , n10442 );
    and g23881 ( n29423 , n28980 , n23091 );
    or g23882 ( n26027 , n2309 , n10591 );
    or g23883 ( n29959 , n22437 , n16343 );
    xnor g23884 ( n5654 , n26563 , n19132 );
    not g23885 ( n17074 , n20345 );
    not g23886 ( n30176 , n9783 );
    not g23887 ( n29727 , n10922 );
    not g23888 ( n6611 , n16393 );
    xnor g23889 ( n2175 , n4513 , n3239 );
    not g23890 ( n14636 , n26052 );
    not g23891 ( n11232 , n15261 );
    or g23892 ( n13588 , n24681 , n18291 );
    nor g23893 ( n29707 , n655 , n21883 );
    nor g23894 ( n31517 , n24794 , n18955 );
    not g23895 ( n28109 , n14268 );
    and g23896 ( n31680 , n7480 , n12930 );
    xnor g23897 ( n4573 , n8359 , n8867 );
    or g23898 ( n18756 , n4105 , n16983 );
    or g23899 ( n27886 , n29668 , n18265 );
    not g23900 ( n16947 , n12208 );
    not g23901 ( n26536 , n7342 );
    not g23902 ( n13432 , n50 );
    nor g23903 ( n31240 , n891 , n22870 );
    or g23904 ( n22648 , n31778 , n29699 );
    not g23905 ( n30578 , n1033 );
    not g23906 ( n25589 , n19680 );
    or g23907 ( n9051 , n8512 , n14817 );
    not g23908 ( n31330 , n8736 );
    not g23909 ( n12893 , n449 );
    not g23910 ( n22420 , n20052 );
    and g23911 ( n12324 , n29798 , n775 );
    not g23912 ( n17001 , n19396 );
    xor g23913 ( n24422 , n7996 , n26998 );
    not g23914 ( n2775 , n7414 );
    nor g23915 ( n27922 , n8773 , n4218 );
    xnor g23916 ( n1260 , n6651 , n3281 );
    and g23917 ( n10275 , n22175 , n26928 );
    and g23918 ( n17222 , n15388 , n15474 );
    not g23919 ( n10316 , n11971 );
    or g23920 ( n8871 , n6987 , n26972 );
    or g23921 ( n15611 , n20158 , n6411 );
    and g23922 ( n12656 , n31251 , n20228 );
    not g23923 ( n24444 , n1229 );
    xnor g23924 ( n29391 , n24000 , n17418 );
    or g23925 ( n19604 , n12750 , n18408 );
    not g23926 ( n28911 , n9939 );
    and g23927 ( n8687 , n13036 , n21779 );
    not g23928 ( n30657 , n16476 );
    xnor g23929 ( n16491 , n2898 , n17305 );
    or g23930 ( n30289 , n8341 , n4055 );
    xnor g23931 ( n14518 , n4908 , n12055 );
    or g23932 ( n28762 , n6527 , n5410 );
    and g23933 ( n13656 , n21390 , n9276 );
    xor g23934 ( n5197 , n7583 , n626 );
    or g23935 ( n22554 , n26944 , n11004 );
    xnor g23936 ( n3942 , n17708 , n27556 );
    not g23937 ( n17148 , n25731 );
    not g23938 ( n13112 , n20895 );
    or g23939 ( n4831 , n18949 , n8271 );
    not g23940 ( n3830 , n6154 );
    not g23941 ( n21520 , n25603 );
    or g23942 ( n23807 , n25556 , n22948 );
    or g23943 ( n975 , n7182 , n7118 );
    or g23944 ( n16066 , n14024 , n6619 );
    xnor g23945 ( n25764 , n789 , n13049 );
    xnor g23946 ( n10305 , n16845 , n1250 );
    xnor g23947 ( n19518 , n2820 , n213 );
    or g23948 ( n16935 , n2400 , n20647 );
    not g23949 ( n29301 , n7930 );
    not g23950 ( n31126 , n30872 );
    xnor g23951 ( n29415 , n19599 , n21137 );
    nor g23952 ( n11316 , n18381 , n16963 );
    or g23953 ( n22359 , n13010 , n29962 );
    or g23954 ( n6488 , n5022 , n14188 );
    or g23955 ( n2342 , n26899 , n2008 );
    or g23956 ( n12134 , n933 , n6611 );
    not g23957 ( n10107 , n7159 );
    and g23958 ( n27009 , n2489 , n9885 );
    not g23959 ( n17010 , n20988 );
    nor g23960 ( n1206 , n5711 , n16655 );
    xnor g23961 ( n21702 , n12121 , n379 );
    not g23962 ( n23596 , n404 );
    nor g23963 ( n28873 , n17766 , n8185 );
    xnor g23964 ( n18369 , n13980 , n7184 );
    or g23965 ( n29461 , n27040 , n6973 );
    xnor g23966 ( n3415 , n14510 , n10682 );
    not g23967 ( n30739 , n7487 );
    nor g23968 ( n23513 , n24531 , n22384 );
    not g23969 ( n6726 , n14160 );
    or g23970 ( n9399 , n30286 , n5671 );
    and g23971 ( n30832 , n17086 , n990 );
    xnor g23972 ( n12012 , n29299 , n27236 );
    xnor g23973 ( n13648 , n15285 , n21448 );
    or g23974 ( n15712 , n549 , n28157 );
    and g23975 ( n5257 , n9510 , n28321 );
    and g23976 ( n17458 , n18818 , n7236 );
    or g23977 ( n10201 , n12180 , n12914 );
    nor g23978 ( n21323 , n8640 , n17966 );
    not g23979 ( n7103 , n28069 );
    or g23980 ( n9194 , n5852 , n10541 );
    or g23981 ( n28928 , n27680 , n15209 );
    not g23982 ( n8166 , n2665 );
    or g23983 ( n5470 , n11375 , n16208 );
    or g23984 ( n5117 , n18041 , n4919 );
    or g23985 ( n25873 , n28776 , n26295 );
    xnor g23986 ( n21758 , n14649 , n14405 );
    not g23987 ( n2488 , n20165 );
    not g23988 ( n6483 , n20960 );
    not g23989 ( n27362 , n24236 );
    not g23990 ( n8655 , n15105 );
    and g23991 ( n18425 , n1534 , n107 );
    and g23992 ( n21061 , n377 , n17160 );
    nor g23993 ( n30888 , n140 , n19244 );
    and g23994 ( n31964 , n31205 , n28022 );
    not g23995 ( n832 , n16968 );
    not g23996 ( n23678 , n2529 );
    xnor g23997 ( n14934 , n14888 , n25213 );
    xnor g23998 ( n4379 , n20489 , n13554 );
    xnor g23999 ( n13266 , n7890 , n14489 );
    not g24000 ( n366 , n11537 );
    not g24001 ( n4499 , n27643 );
    or g24002 ( n2390 , n25708 , n6983 );
    or g24003 ( n16768 , n24963 , n13904 );
    not g24004 ( n2997 , n9376 );
    and g24005 ( n9006 , n2194 , n16482 );
    nor g24006 ( n6208 , n20656 , n27419 );
    nor g24007 ( n2616 , n7209 , n291 );
    not g24008 ( n23061 , n17886 );
    not g24009 ( n21452 , n97 );
    or g24010 ( n6759 , n25927 , n4233 );
    or g24011 ( n11939 , n1972 , n5512 );
    not g24012 ( n9059 , n22123 );
    or g24013 ( n29613 , n24145 , n27495 );
    or g24014 ( n27138 , n31284 , n18186 );
    not g24015 ( n23823 , n27724 );
    xnor g24016 ( n18793 , n2082 , n14669 );
    not g24017 ( n27881 , n6720 );
    xnor g24018 ( n27414 , n24132 , n256 );
    xnor g24019 ( n24987 , n365 , n5949 );
    xnor g24020 ( n3557 , n552 , n30423 );
    or g24021 ( n31929 , n20781 , n13875 );
    xnor g24022 ( n10620 , n4559 , n15057 );
    or g24023 ( n8156 , n27649 , n9126 );
    or g24024 ( n11831 , n21111 , n6325 );
    xnor g24025 ( n15460 , n25905 , n5493 );
    or g24026 ( n371 , n15320 , n25204 );
    or g24027 ( n21538 , n14202 , n13370 );
    not g24028 ( n8398 , n20861 );
    not g24029 ( n16213 , n28204 );
    or g24030 ( n24825 , n26412 , n27246 );
    not g24031 ( n22095 , n21463 );
    and g24032 ( n2111 , n3801 , n10758 );
    not g24033 ( n12496 , n22287 );
    not g24034 ( n23715 , n6207 );
    not g24035 ( n30233 , n16953 );
    or g24036 ( n26921 , n29422 , n21634 );
    or g24037 ( n20725 , n1044 , n6260 );
    nor g24038 ( n6975 , n15935 , n18085 );
    xnor g24039 ( n30282 , n21035 , n13695 );
    not g24040 ( n25938 , n7098 );
    not g24041 ( n6787 , n5948 );
    not g24042 ( n2620 , n16441 );
    or g24043 ( n12603 , n15600 , n24208 );
    xnor g24044 ( n20164 , n10384 , n22180 );
    or g24045 ( n14972 , n30464 , n27718 );
    not g24046 ( n15527 , n13759 );
    nor g24047 ( n27466 , n5900 , n23196 );
    or g24048 ( n27596 , n10018 , n17483 );
    not g24049 ( n25028 , n925 );
    not g24050 ( n14464 , n11063 );
    not g24051 ( n10310 , n19433 );
    or g24052 ( n845 , n2694 , n28170 );
    not g24053 ( n28718 , n13266 );
    or g24054 ( n28855 , n20177 , n23099 );
    not g24055 ( n646 , n15795 );
    or g24056 ( n6235 , n8919 , n28913 );
    or g24057 ( n17708 , n13082 , n24277 );
    xnor g24058 ( n3795 , n12915 , n1265 );
    xnor g24059 ( n10136 , n9294 , n1686 );
    nor g24060 ( n17362 , n2963 , n25260 );
    xnor g24061 ( n2848 , n652 , n30108 );
    xnor g24062 ( n7482 , n25711 , n14178 );
    not g24063 ( n23511 , n4529 );
    xnor g24064 ( n17489 , n3936 , n21188 );
    xnor g24065 ( n2556 , n8986 , n5313 );
    or g24066 ( n19178 , n16075 , n8524 );
    not g24067 ( n12286 , n20649 );
    nor g24068 ( n23364 , n20168 , n12688 );
    nor g24069 ( n8012 , n20582 , n30410 );
    not g24070 ( n20420 , n20771 );
    nor g24071 ( n770 , n2665 , n26866 );
    or g24072 ( n11848 , n29998 , n16660 );
    nor g24073 ( n15502 , n29444 , n7844 );
    nor g24074 ( n26097 , n20796 , n19886 );
    nor g24075 ( n70 , n1086 , n21973 );
    or g24076 ( n18066 , n13134 , n3125 );
    or g24077 ( n22282 , n19097 , n2043 );
    or g24078 ( n22353 , n17997 , n25044 );
    xnor g24079 ( n19926 , n28296 , n18861 );
    not g24080 ( n30964 , n30259 );
    not g24081 ( n30126 , n10067 );
    xnor g24082 ( n18880 , n14660 , n4339 );
    and g24083 ( n24992 , n31771 , n19447 );
    and g24084 ( n17121 , n29644 , n28056 );
    nor g24085 ( n30097 , n12446 , n1216 );
    or g24086 ( n14309 , n25236 , n10604 );
    xnor g24087 ( n3443 , n28889 , n30974 );
    not g24088 ( n23820 , n31424 );
    or g24089 ( n1222 , n13529 , n1061 );
    xnor g24090 ( n8112 , n13789 , n7407 );
    and g24091 ( n26278 , n9560 , n18535 );
    xnor g24092 ( n24363 , n23048 , n12831 );
    or g24093 ( n11926 , n23891 , n11709 );
    nor g24094 ( n14616 , n1635 , n2296 );
    not g24095 ( n2431 , n17530 );
    not g24096 ( n22924 , n28634 );
    and g24097 ( n24813 , n19795 , n4353 );
    or g24098 ( n17816 , n24828 , n9551 );
    and g24099 ( n4320 , n17088 , n24941 );
    or g24100 ( n22720 , n28496 , n8895 );
    nor g24101 ( n30569 , n14039 , n10627 );
    xnor g24102 ( n11494 , n10780 , n26974 );
    and g24103 ( n20584 , n2689 , n11300 );
    not g24104 ( n13148 , n22793 );
    xnor g24105 ( n17929 , n1856 , n20390 );
    xnor g24106 ( n4982 , n24097 , n17675 );
    xnor g24107 ( n14311 , n24250 , n27474 );
    or g24108 ( n24098 , n22807 , n14786 );
    xnor g24109 ( n8849 , n14670 , n14962 );
    not g24110 ( n11573 , n8919 );
    not g24111 ( n20167 , n4247 );
    and g24112 ( n20502 , n13603 , n7959 );
    or g24113 ( n5010 , n12035 , n2712 );
    not g24114 ( n18761 , n17811 );
    xnor g24115 ( n20194 , n17775 , n22104 );
    xnor g24116 ( n13969 , n20441 , n31545 );
    nor g24117 ( n16673 , n11866 , n31500 );
    or g24118 ( n26759 , n27591 , n29746 );
    nor g24119 ( n2667 , n6319 , n31141 );
    xnor g24120 ( n12638 , n28045 , n21154 );
    or g24121 ( n25465 , n31840 , n3402 );
    not g24122 ( n9734 , n26798 );
    and g24123 ( n13 , n31742 , n11715 );
    not g24124 ( n236 , n24899 );
    or g24125 ( n18994 , n8003 , n6607 );
    nor g24126 ( n1759 , n594 , n16560 );
    xnor g24127 ( n1258 , n5217 , n7133 );
    xnor g24128 ( n24817 , n722 , n9717 );
    and g24129 ( n6589 , n11114 , n25009 );
    not g24130 ( n20975 , n16000 );
    not g24131 ( n27199 , n12275 );
    xnor g24132 ( n16345 , n693 , n21942 );
    nor g24133 ( n2832 , n11152 , n5279 );
    or g24134 ( n13042 , n29681 , n27769 );
    xnor g24135 ( n29806 , n3822 , n3688 );
    xnor g24136 ( n29711 , n21516 , n13672 );
    or g24137 ( n13769 , n33 , n19590 );
    xnor g24138 ( n16711 , n4464 , n30404 );
    xnor g24139 ( n19556 , n28356 , n3312 );
    not g24140 ( n23856 , n27866 );
    xnor g24141 ( n18981 , n16873 , n20181 );
    xnor g24142 ( n10865 , n6062 , n12260 );
    and g24143 ( n24436 , n8772 , n28290 );
    xor g24144 ( n6394 , n13733 , n2551 );
    nor g24145 ( n12916 , n13980 , n15204 );
    or g24146 ( n9131 , n28542 , n29873 );
    xnor g24147 ( n9362 , n2710 , n30814 );
    or g24148 ( n2463 , n1648 , n28601 );
    not g24149 ( n10427 , n13726 );
    not g24150 ( n15081 , n17745 );
    nor g24151 ( n30591 , n19279 , n21875 );
    or g24152 ( n27664 , n911 , n15789 );
    xnor g24153 ( n3113 , n23263 , n8083 );
    and g24154 ( n27255 , n5730 , n19537 );
    xnor g24155 ( n3070 , n2052 , n18230 );
    not g24156 ( n25233 , n8451 );
    not g24157 ( n24589 , n27475 );
    xor g24158 ( n24358 , n7329 , n2330 );
    or g24159 ( n30143 , n26275 , n24059 );
    and g24160 ( n17232 , n21331 , n23600 );
    xnor g24161 ( n16882 , n18732 , n3156 );
    and g24162 ( n10293 , n10717 , n25515 );
    or g24163 ( n27042 , n27408 , n439 );
    or g24164 ( n24885 , n1765 , n2488 );
    not g24165 ( n8969 , n8151 );
    not g24166 ( n21275 , n25026 );
    and g24167 ( n1813 , n22073 , n6643 );
    or g24168 ( n24395 , n30691 , n9820 );
    or g24169 ( n4677 , n12298 , n11506 );
    not g24170 ( n17432 , n11287 );
    nor g24171 ( n17616 , n21817 , n821 );
    and g24172 ( n8050 , n13055 , n28214 );
    or g24173 ( n7373 , n27311 , n17268 );
    xnor g24174 ( n4495 , n4742 , n8445 );
    not g24175 ( n23283 , n4003 );
    and g24176 ( n10272 , n20077 , n14628 );
    or g24177 ( n5333 , n31202 , n13388 );
    xnor g24178 ( n828 , n321 , n7264 );
    xnor g24179 ( n18235 , n31281 , n13895 );
    xnor g24180 ( n13811 , n27100 , n22623 );
    nor g24181 ( n18946 , n19962 , n31308 );
    xnor g24182 ( n28337 , n14815 , n17466 );
    not g24183 ( n23595 , n19814 );
    buf g24184 ( n8931 , n11981 );
    xnor g24185 ( n24236 , n18031 , n20759 );
    not g24186 ( n24857 , n2490 );
    not g24187 ( n27966 , n31739 );
    or g24188 ( n6101 , n14290 , n1100 );
    xnor g24189 ( n10608 , n23766 , n19118 );
    not g24190 ( n607 , n15035 );
    not g24191 ( n28705 , n31986 );
    or g24192 ( n14353 , n7028 , n8144 );
    not g24193 ( n18419 , n1031 );
    xnor g24194 ( n21989 , n6186 , n26228 );
    not g24195 ( n10049 , n21204 );
    nor g24196 ( n18713 , n22788 , n11056 );
    or g24197 ( n31674 , n22298 , n27079 );
    xnor g24198 ( n10101 , n6415 , n22451 );
    and g24199 ( n13542 , n29090 , n23040 );
    nor g24200 ( n24985 , n2483 , n18955 );
    or g24201 ( n21811 , n29904 , n12723 );
    or g24202 ( n21368 , n13613 , n1860 );
    or g24203 ( n6877 , n18356 , n29590 );
    or g24204 ( n8362 , n23720 , n29761 );
    xnor g24205 ( n13932 , n13909 , n14148 );
    or g24206 ( n3900 , n12109 , n13828 );
    or g24207 ( n27222 , n26788 , n1772 );
    not g24208 ( n4494 , n27429 );
    xnor g24209 ( n19283 , n17889 , n25095 );
    or g24210 ( n17975 , n29236 , n17968 );
    not g24211 ( n31694 , n10123 );
    nor g24212 ( n13031 , n6849 , n27381 );
    not g24213 ( n31214 , n22142 );
    xor g24214 ( n31887 , n9790 , n18870 );
    not g24215 ( n16842 , n7354 );
    or g24216 ( n20835 , n14549 , n21946 );
    or g24217 ( n30885 , n6655 , n23597 );
    xnor g24218 ( n8483 , n22652 , n20960 );
    or g24219 ( n4053 , n2966 , n370 );
    xnor g24220 ( n23293 , n13874 , n1546 );
    not g24221 ( n19830 , n12080 );
    and g24222 ( n1610 , n6679 , n803 );
    not g24223 ( n9669 , n29015 );
    or g24224 ( n13000 , n22692 , n8424 );
    and g24225 ( n25352 , n23945 , n30661 );
    or g24226 ( n23851 , n29165 , n5724 );
    xnor g24227 ( n18683 , n5758 , n5270 );
    xnor g24228 ( n22829 , n12848 , n22828 );
    not g24229 ( n16134 , n21597 );
    or g24230 ( n1237 , n18553 , n19703 );
    and g24231 ( n19276 , n6572 , n4400 );
    not g24232 ( n12045 , n18977 );
    not g24233 ( n3574 , n17093 );
    not g24234 ( n6885 , n1348 );
    or g24235 ( n11495 , n2777 , n21137 );
    or g24236 ( n16510 , n19221 , n1131 );
    or g24237 ( n9597 , n1540 , n25111 );
    or g24238 ( n9817 , n30829 , n18748 );
    or g24239 ( n7223 , n8183 , n14419 );
    nor g24240 ( n22486 , n1423 , n32017 );
    not g24241 ( n13420 , n9884 );
    or g24242 ( n7238 , n2370 , n23967 );
    nor g24243 ( n24333 , n20012 , n13688 );
    xnor g24244 ( n7896 , n20163 , n1007 );
    nor g24245 ( n2207 , n4374 , n21553 );
    not g24246 ( n10043 , n29895 );
    not g24247 ( n12526 , n20982 );
    xnor g24248 ( n16468 , n31273 , n30472 );
    not g24249 ( n14036 , n1830 );
    not g24250 ( n20028 , n25993 );
    not g24251 ( n31849 , n4335 );
    nor g24252 ( n13160 , n22529 , n31257 );
    nor g24253 ( n26026 , n4649 , n10518 );
    and g24254 ( n18287 , n29017 , n27523 );
    not g24255 ( n29378 , n13382 );
    or g24256 ( n6665 , n20286 , n14600 );
    not g24257 ( n17743 , n7473 );
    xnor g24258 ( n252 , n22802 , n31722 );
    xnor g24259 ( n265 , n23483 , n4335 );
    xnor g24260 ( n6928 , n16960 , n78 );
    nor g24261 ( n22425 , n11736 , n20463 );
    nor g24262 ( n2234 , n14503 , n19357 );
    xnor g24263 ( n11485 , n8021 , n5517 );
    or g24264 ( n22078 , n8717 , n17940 );
    and g24265 ( n25083 , n23657 , n23681 );
    not g24266 ( n7208 , n8462 );
    or g24267 ( n15072 , n23728 , n5217 );
    or g24268 ( n8786 , n19862 , n900 );
    not g24269 ( n22227 , n25202 );
    not g24270 ( n17002 , n30018 );
    xnor g24271 ( n13074 , n9835 , n26004 );
    or g24272 ( n16596 , n27717 , n20477 );
    not g24273 ( n13496 , n23934 );
    not g24274 ( n29560 , n8864 );
    or g24275 ( n1436 , n21984 , n8318 );
    and g24276 ( n17735 , n7756 , n25328 );
    not g24277 ( n2762 , n19021 );
    not g24278 ( n2589 , n22937 );
    and g24279 ( n29701 , n26000 , n26779 );
    and g24280 ( n25375 , n6289 , n21825 );
    or g24281 ( n13699 , n3292 , n31859 );
    nor g24282 ( n4306 , n205 , n28575 );
    not g24283 ( n3753 , n14239 );
    or g24284 ( n3629 , n19922 , n221 );
    xnor g24285 ( n13711 , n24253 , n25813 );
    or g24286 ( n8703 , n15427 , n31646 );
    not g24287 ( n3486 , n20968 );
    or g24288 ( n2944 , n24721 , n2641 );
    and g24289 ( n14210 , n30147 , n13294 );
    not g24290 ( n17774 , n21136 );
    not g24291 ( n24881 , n17798 );
    and g24292 ( n13636 , n23609 , n2662 );
    not g24293 ( n26640 , n30199 );
    not g24294 ( n27019 , n9956 );
    nor g24295 ( n27375 , n4111 , n16891 );
    xnor g24296 ( n25135 , n19031 , n25438 );
    not g24297 ( n2845 , n2368 );
    xnor g24298 ( n31153 , n1648 , n9718 );
    nor g24299 ( n16568 , n10772 , n8514 );
    nor g24300 ( n22838 , n10847 , n19292 );
    not g24301 ( n14468 , n4318 );
    not g24302 ( n22193 , n16241 );
    or g24303 ( n27159 , n18778 , n15160 );
    and g24304 ( n3389 , n14524 , n6551 );
    or g24305 ( n15630 , n9374 , n1722 );
    and g24306 ( n16513 , n28764 , n12844 );
    xnor g24307 ( n3991 , n16416 , n8849 );
    xnor g24308 ( n13090 , n19537 , n17952 );
    nor g24309 ( n18434 , n17840 , n1054 );
    xnor g24310 ( n12320 , n28198 , n25470 );
    xnor g24311 ( n15891 , n11865 , n19712 );
    and g24312 ( n5216 , n25990 , n30307 );
    or g24313 ( n19993 , n29424 , n30651 );
    buf g24314 ( n2301 , n30336 );
    nor g24315 ( n1790 , n18389 , n25497 );
    and g24316 ( n28602 , n24215 , n2172 );
    or g24317 ( n992 , n13241 , n25394 );
    xnor g24318 ( n10417 , n18592 , n18726 );
    and g24319 ( n8952 , n1591 , n20836 );
    xnor g24320 ( n11778 , n1044 , n18329 );
    xnor g24321 ( n14761 , n15972 , n28338 );
    xor g24322 ( n4934 , n5556 , n25489 );
    or g24323 ( n15865 , n16557 , n13371 );
    xnor g24324 ( n19194 , n640 , n11059 );
    xnor g24325 ( n10416 , n6662 , n10490 );
    and g24326 ( n7865 , n13386 , n57 );
    nor g24327 ( n6467 , n3822 , n23097 );
    xnor g24328 ( n30162 , n30630 , n23499 );
    or g24329 ( n3503 , n25533 , n16327 );
    xnor g24330 ( n19793 , n24446 , n22440 );
    and g24331 ( n5353 , n8691 , n8690 );
    not g24332 ( n31513 , n10555 );
    and g24333 ( n30191 , n16590 , n15841 );
    not g24334 ( n4793 , n12061 );
    not g24335 ( n23133 , n10261 );
    or g24336 ( n17114 , n29044 , n10661 );
    not g24337 ( n28463 , n25514 );
    and g24338 ( n19541 , n1189 , n27257 );
    and g24339 ( n2531 , n3544 , n6388 );
    xnor g24340 ( n27530 , n2627 , n4918 );
    and g24341 ( n4212 , n16501 , n18368 );
    or g24342 ( n11696 , n23943 , n4768 );
    or g24343 ( n3742 , n21395 , n23845 );
    not g24344 ( n18895 , n19594 );
    or g24345 ( n4603 , n15396 , n2731 );
    not g24346 ( n4305 , n7880 );
    xor g24347 ( n29195 , n14878 , n24834 );
    xor g24348 ( n26261 , n31734 , n19035 );
    or g24349 ( n11303 , n3765 , n7915 );
    nor g24350 ( n10227 , n6888 , n6674 );
    not g24351 ( n17622 , n9500 );
    xnor g24352 ( n14288 , n31593 , n15371 );
    and g24353 ( n15599 , n25155 , n27744 );
    or g24354 ( n15801 , n5354 , n22566 );
    not g24355 ( n3233 , n5420 );
    not g24356 ( n9721 , n19614 );
    or g24357 ( n21074 , n20373 , n1140 );
    xnor g24358 ( n4315 , n13387 , n14925 );
    or g24359 ( n9089 , n3820 , n6026 );
    not g24360 ( n18901 , n6760 );
    or g24361 ( n16886 , n6376 , n4721 );
    or g24362 ( n6265 , n10619 , n26284 );
    and g24363 ( n30891 , n10342 , n9032 );
    or g24364 ( n19119 , n22075 , n26624 );
    xnor g24365 ( n8 , n19700 , n30003 );
    xnor g24366 ( n16643 , n30218 , n18612 );
    or g24367 ( n14433 , n24077 , n17360 );
    xnor g24368 ( n2876 , n24211 , n10775 );
    xnor g24369 ( n15806 , n21996 , n3436 );
    and g24370 ( n7057 , n5726 , n15465 );
    xnor g24371 ( n22381 , n18569 , n2047 );
    xnor g24372 ( n1848 , n3041 , n1467 );
    not g24373 ( n29243 , n29114 );
    nor g24374 ( n12697 , n29668 , n24415 );
    and g24375 ( n24135 , n9231 , n8500 );
    and g24376 ( n19917 , n8021 , n11230 );
    not g24377 ( n27001 , n1037 );
    or g24378 ( n29405 , n18259 , n24258 );
    xnor g24379 ( n12356 , n22845 , n1670 );
    not g24380 ( n6491 , n20350 );
    xnor g24381 ( n31815 , n29090 , n20799 );
    buf g24382 ( n9134 , n21282 );
    or g24383 ( n14113 , n107 , n15348 );
    nor g24384 ( n30840 , n12478 , n16019 );
    and g24385 ( n18748 , n18721 , n31636 );
    and g24386 ( n30400 , n6665 , n31527 );
    and g24387 ( n13311 , n19608 , n30847 );
    or g24388 ( n29601 , n20336 , n13885 );
    xnor g24389 ( n5252 , n8978 , n13200 );
    not g24390 ( n6283 , n27266 );
    not g24391 ( n22567 , n11264 );
    or g24392 ( n30510 , n26737 , n11586 );
    not g24393 ( n5290 , n17609 );
    and g24394 ( n25962 , n7608 , n16638 );
    and g24395 ( n28699 , n16511 , n28444 );
    and g24396 ( n13302 , n17513 , n15659 );
    xnor g24397 ( n28520 , n10477 , n2883 );
    nor g24398 ( n23906 , n16658 , n13351 );
    and g24399 ( n10661 , n30294 , n14251 );
    xnor g24400 ( n27086 , n7792 , n9555 );
    nor g24401 ( n20941 , n21288 , n11929 );
    xnor g24402 ( n17390 , n30002 , n29471 );
    or g24403 ( n26697 , n9290 , n18458 );
    not g24404 ( n17459 , n26774 );
    not g24405 ( n21553 , n2027 );
    not g24406 ( n17580 , n7626 );
    or g24407 ( n20564 , n28444 , n16511 );
    and g24408 ( n8247 , n4726 , n18277 );
    and g24409 ( n26648 , n19674 , n3644 );
    or g24410 ( n8121 , n1847 , n4473 );
    nor g24411 ( n30068 , n3166 , n15718 );
    nor g24412 ( n19910 , n10805 , n9674 );
    not g24413 ( n31110 , n471 );
    xnor g24414 ( n19021 , n3374 , n14966 );
    and g24415 ( n4876 , n3373 , n7816 );
    and g24416 ( n24907 , n0 , n480 );
    xnor g24417 ( n3726 , n21238 , n29744 );
    nor g24418 ( n19369 , n554 , n5251 );
    not g24419 ( n12879 , n10158 );
    and g24420 ( n15196 , n3627 , n25592 );
    not g24421 ( n6163 , n2971 );
    and g24422 ( n20389 , n5063 , n15326 );
    not g24423 ( n3566 , n28179 );
    xnor g24424 ( n22125 , n23509 , n17452 );
    xnor g24425 ( n28661 , n9011 , n20198 );
    or g24426 ( n4955 , n11072 , n9790 );
    and g24427 ( n26187 , n15999 , n23097 );
    xnor g24428 ( n21588 , n6052 , n3214 );
    not g24429 ( n20788 , n25192 );
    and g24430 ( n8785 , n22265 , n31547 );
    and g24431 ( n25404 , n7167 , n24859 );
    xnor g24432 ( n11289 , n5863 , n9322 );
    nor g24433 ( n26106 , n16274 , n16561 );
    xnor g24434 ( n17863 , n16395 , n31661 );
    not g24435 ( n13580 , n27501 );
    xnor g24436 ( n18303 , n4303 , n22469 );
    buf g24437 ( n20052 , n22236 );
    not g24438 ( n25743 , n25629 );
    not g24439 ( n13796 , n21513 );
    xnor g24440 ( n14753 , n5156 , n921 );
    xnor g24441 ( n10445 , n31108 , n3289 );
    nor g24442 ( n25457 , n24358 , n14527 );
    not g24443 ( n3453 , n16345 );
    xnor g24444 ( n16393 , n7327 , n20346 );
    xnor g24445 ( n6310 , n27270 , n30106 );
    not g24446 ( n31306 , n8477 );
    xnor g24447 ( n14868 , n471 , n6223 );
    or g24448 ( n28966 , n21926 , n11506 );
    xnor g24449 ( n18897 , n4827 , n12677 );
    or g24450 ( n17009 , n1497 , n1950 );
    not g24451 ( n442 , n5160 );
    not g24452 ( n16276 , n12963 );
    not g24453 ( n28580 , n10467 );
    xnor g24454 ( n15026 , n21713 , n22093 );
    xnor g24455 ( n9605 , n2180 , n6527 );
    and g24456 ( n9688 , n20654 , n8033 );
    xnor g24457 ( n28115 , n26052 , n27077 );
    and g24458 ( n6520 , n15423 , n17800 );
    or g24459 ( n4885 , n17421 , n4180 );
    xnor g24460 ( n18508 , n28231 , n19396 );
    or g24461 ( n9158 , n24325 , n16086 );
    or g24462 ( n22812 , n15955 , n902 );
    not g24463 ( n26429 , n14197 );
    or g24464 ( n8587 , n4399 , n10330 );
    xnor g24465 ( n17657 , n21190 , n7551 );
    xnor g24466 ( n30776 , n4312 , n1897 );
    nor g24467 ( n31229 , n4194 , n19295 );
    xnor g24468 ( n14780 , n5473 , n3641 );
    or g24469 ( n27458 , n23488 , n7574 );
    not g24470 ( n13376 , n18831 );
    or g24471 ( n17811 , n20495 , n4470 );
    not g24472 ( n16112 , n21383 );
    not g24473 ( n10047 , n5747 );
    xnor g24474 ( n10800 , n22321 , n18153 );
    or g24475 ( n9030 , n5028 , n26763 );
    or g24476 ( n29605 , n6957 , n18284 );
    and g24477 ( n22314 , n7548 , n2665 );
    xnor g24478 ( n25877 , n21881 , n32016 );
    or g24479 ( n27349 , n23577 , n30461 );
    or g24480 ( n15546 , n29989 , n27061 );
    not g24481 ( n26387 , n5400 );
    not g24482 ( n13034 , n2741 );
    or g24483 ( n5263 , n27339 , n21795 );
    not g24484 ( n6615 , n24201 );
    nor g24485 ( n1804 , n18883 , n8665 );
    xnor g24486 ( n31639 , n4513 , n24907 );
    and g24487 ( n31081 , n22822 , n26703 );
    xnor g24488 ( n3596 , n28446 , n17415 );
    not g24489 ( n20120 , n29042 );
    or g24490 ( n23031 , n28548 , n6975 );
    or g24491 ( n8517 , n14728 , n6746 );
    and g24492 ( n18179 , n10545 , n9516 );
    not g24493 ( n16259 , n8433 );
    buf g24494 ( n31338 , n17790 );
    xnor g24495 ( n30803 , n29569 , n16113 );
    nor g24496 ( n21184 , n5126 , n7438 );
    or g24497 ( n29706 , n22015 , n31900 );
    xnor g24498 ( n21570 , n1949 , n26939 );
    not g24499 ( n22021 , n30622 );
    not g24500 ( n8355 , n32024 );
    and g24501 ( n2926 , n25131 , n11695 );
    xnor g24502 ( n25895 , n3536 , n26505 );
    or g24503 ( n22445 , n30112 , n5405 );
    nor g24504 ( n15952 , n21122 , n7655 );
    and g24505 ( n270 , n16997 , n8988 );
    and g24506 ( n20855 , n2671 , n17275 );
    or g24507 ( n11180 , n25276 , n4844 );
    and g24508 ( n27924 , n18574 , n32013 );
    or g24509 ( n3841 , n26244 , n23616 );
    or g24510 ( n30630 , n4600 , n21922 );
    not g24511 ( n10183 , n5432 );
    xnor g24512 ( n19775 , n13129 , n17051 );
    and g24513 ( n28693 , n5023 , n25293 );
    or g24514 ( n23307 , n8171 , n25045 );
    not g24515 ( n24158 , n28712 );
    or g24516 ( n28784 , n9447 , n25523 );
    and g24517 ( n30403 , n5199 , n17128 );
    or g24518 ( n1472 , n893 , n28393 );
    or g24519 ( n23935 , n14538 , n1567 );
    and g24520 ( n20682 , n27726 , n8372 );
    not g24521 ( n17008 , n23788 );
    xnor g24522 ( n21980 , n1703 , n20168 );
    not g24523 ( n9763 , n10537 );
    not g24524 ( n3138 , n18980 );
    and g24525 ( n12914 , n1911 , n3391 );
    not g24526 ( n17334 , n15362 );
    or g24527 ( n27838 , n28667 , n2841 );
    or g24528 ( n4353 , n18104 , n7384 );
    not g24529 ( n8544 , n25756 );
    xnor g24530 ( n15007 , n19377 , n8153 );
    not g24531 ( n4688 , n6128 );
    and g24532 ( n12288 , n14238 , n27276 );
    and g24533 ( n26842 , n10828 , n864 );
    and g24534 ( n16641 , n2672 , n7135 );
    not g24535 ( n18656 , n19294 );
    not g24536 ( n13756 , n21880 );
    and g24537 ( n4109 , n27055 , n31281 );
    nor g24538 ( n24711 , n11361 , n13172 );
    not g24539 ( n1871 , n16113 );
    or g24540 ( n4406 , n2954 , n9576 );
    or g24541 ( n19225 , n14374 , n17292 );
    buf g24542 ( n26109 , n12338 );
    or g24543 ( n6490 , n10864 , n18062 );
    and g24544 ( n22843 , n2519 , n16710 );
    nor g24545 ( n17911 , n20825 , n12011 );
    xnor g24546 ( n10446 , n18064 , n17336 );
    not g24547 ( n5205 , n2235 );
    or g24548 ( n18353 , n18271 , n28348 );
    not g24549 ( n18511 , n3873 );
    or g24550 ( n7213 , n15016 , n2015 );
    not g24551 ( n22441 , n25201 );
    not g24552 ( n25649 , n17798 );
    xnor g24553 ( n26918 , n2731 , n24377 );
    xnor g24554 ( n17718 , n27317 , n26758 );
    nor g24555 ( n415 , n20746 , n29043 );
    not g24556 ( n13307 , n20996 );
    and g24557 ( n11929 , n27119 , n3127 );
    or g24558 ( n7602 , n15432 , n765 );
    not g24559 ( n14027 , n12143 );
    xnor g24560 ( n24747 , n30887 , n10034 );
    not g24561 ( n8776 , n8355 );
    not g24562 ( n30427 , n6266 );
    xnor g24563 ( n10649 , n31754 , n23620 );
    or g24564 ( n133 , n11727 , n23573 );
    not g24565 ( n10913 , n8510 );
    or g24566 ( n13719 , n3659 , n11985 );
    not g24567 ( n28243 , n24698 );
    not g24568 ( n19493 , n14542 );
    not g24569 ( n26580 , n4935 );
    xnor g24570 ( n28960 , n15814 , n9703 );
    xnor g24571 ( n27075 , n26406 , n29569 );
    xnor g24572 ( n27022 , n7937 , n7749 );
    not g24573 ( n20005 , n18164 );
    or g24574 ( n9476 , n5313 , n12757 );
    and g24575 ( n12225 , n16939 , n24076 );
    or g24576 ( n18299 , n18483 , n288 );
    xor g24577 ( n23100 , n10046 , n19239 );
    nor g24578 ( n8738 , n6995 , n27439 );
    or g24579 ( n4269 , n1385 , n9735 );
    and g24580 ( n14090 , n17774 , n28084 );
    or g24581 ( n19875 , n28844 , n6000 );
    and g24582 ( n10683 , n19326 , n27034 );
    xnor g24583 ( n26017 , n5910 , n11477 );
    xnor g24584 ( n19769 , n28624 , n23111 );
    xnor g24585 ( n25382 , n5150 , n5873 );
    not g24586 ( n17030 , n26708 );
    xor g24587 ( n28523 , n773 , n25753 );
    xnor g24588 ( n20721 , n23652 , n27995 );
    not g24589 ( n1648 , n18208 );
    xnor g24590 ( n1901 , n12949 , n20433 );
    xnor g24591 ( n22138 , n18709 , n23060 );
    or g24592 ( n5225 , n13647 , n17353 );
    xor g24593 ( n19642 , n1674 , n3176 );
    not g24594 ( n10395 , n13057 );
    or g24595 ( n26063 , n20155 , n14624 );
    not g24596 ( n17765 , n19879 );
    and g24597 ( n5810 , n9874 , n262 );
    nor g24598 ( n20045 , n24213 , n2821 );
    or g24599 ( n31726 , n30080 , n4937 );
    xnor g24600 ( n22730 , n1704 , n26929 );
    or g24601 ( n12281 , n9154 , n6124 );
    and g24602 ( n23825 , n7646 , n15698 );
    and g24603 ( n25907 , n19968 , n544 );
    and g24604 ( n14417 , n14252 , n29665 );
    or g24605 ( n22 , n30220 , n18854 );
    not g24606 ( n10357 , n31379 );
    not g24607 ( n22296 , n2347 );
    not g24608 ( n28310 , n29065 );
    xnor g24609 ( n27295 , n9501 , n9624 );
    or g24610 ( n377 , n19150 , n13928 );
    and g24611 ( n1466 , n20277 , n31632 );
    or g24612 ( n12735 , n6238 , n16120 );
    or g24613 ( n28316 , n6916 , n31571 );
    xnor g24614 ( n12623 , n21085 , n621 );
    xnor g24615 ( n20270 , n22483 , n16205 );
    and g24616 ( n14949 , n3484 , n24377 );
    buf g24617 ( n11169 , n7818 );
    or g24618 ( n9658 , n6481 , n12341 );
    and g24619 ( n4998 , n28508 , n2743 );
    or g24620 ( n20173 , n4799 , n9721 );
    or g24621 ( n16919 , n29571 , n31867 );
    and g24622 ( n27419 , n31936 , n15284 );
    nor g24623 ( n19259 , n24443 , n25148 );
    xnor g24624 ( n31077 , n16668 , n18235 );
    or g24625 ( n27950 , n3463 , n19332 );
    and g24626 ( n9745 , n11773 , n3366 );
    xnor g24627 ( n9377 , n31633 , n10451 );
    xnor g24628 ( n6739 , n14126 , n7847 );
    or g24629 ( n5762 , n25758 , n21345 );
    not g24630 ( n25066 , n10905 );
    or g24631 ( n26965 , n26455 , n25266 );
    or g24632 ( n6264 , n2644 , n31969 );
    not g24633 ( n19122 , n14504 );
    nor g24634 ( n28483 , n27901 , n28269 );
    xor g24635 ( n7400 , n16964 , n11367 );
    not g24636 ( n5208 , n9769 );
    xnor g24637 ( n22716 , n31705 , n2459 );
    nor g24638 ( n17697 , n8244 , n16445 );
    not g24639 ( n23487 , n24583 );
    not g24640 ( n21 , n12465 );
    xor g24641 ( n20864 , n645 , n31727 );
    xnor g24642 ( n26378 , n2115 , n3133 );
    or g24643 ( n21554 , n4740 , n14532 );
    xnor g24644 ( n8397 , n4206 , n9310 );
    or g24645 ( n9663 , n763 , n14361 );
    or g24646 ( n8976 , n15776 , n11048 );
    and g24647 ( n8857 , n19818 , n12992 );
    xnor g24648 ( n10304 , n26598 , n11060 );
    or g24649 ( n23682 , n1290 , n7164 );
    or g24650 ( n2151 , n2951 , n14737 );
    or g24651 ( n1263 , n20495 , n30525 );
    or g24652 ( n3304 , n13146 , n28814 );
    not g24653 ( n31828 , n4201 );
    and g24654 ( n15786 , n29312 , n2907 );
    nor g24655 ( n12520 , n27093 , n5566 );
    xnor g24656 ( n11411 , n15346 , n15939 );
    or g24657 ( n29136 , n4404 , n11729 );
    or g24658 ( n2456 , n1400 , n4852 );
    and g24659 ( n17825 , n2750 , n88 );
    not g24660 ( n30720 , n30019 );
    not g24661 ( n20398 , n21778 );
    xnor g24662 ( n513 , n26198 , n5759 );
    or g24663 ( n7237 , n15098 , n21048 );
    not g24664 ( n13706 , n21070 );
    xnor g24665 ( n1602 , n22441 , n19299 );
    and g24666 ( n27014 , n26437 , n29302 );
    and g24667 ( n22948 , n11173 , n3617 );
    and g24668 ( n31363 , n11163 , n12332 );
    not g24669 ( n29643 , n20332 );
    and g24670 ( n17056 , n1673 , n24879 );
    not g24671 ( n21786 , n27783 );
    or g24672 ( n5874 , n4657 , n24169 );
    not g24673 ( n6016 , n19808 );
    and g24674 ( n24239 , n3946 , n1107 );
    and g24675 ( n30990 , n12089 , n21285 );
    and g24676 ( n2124 , n18480 , n4855 );
    and g24677 ( n21238 , n28253 , n2501 );
    xor g24678 ( n23246 , n28855 , n14106 );
    or g24679 ( n16693 , n26647 , n3233 );
    xor g24680 ( n13661 , n17070 , n20205 );
    or g24681 ( n20758 , n22076 , n29750 );
    or g24682 ( n2028 , n6246 , n4033 );
    xnor g24683 ( n23464 , n23328 , n6454 );
    and g24684 ( n5478 , n29128 , n29127 );
    xnor g24685 ( n12535 , n19880 , n775 );
    xnor g24686 ( n28475 , n26224 , n17497 );
    xor g24687 ( n19770 , n13592 , n24812 );
    not g24688 ( n4594 , n18181 );
    and g24689 ( n13718 , n24433 , n21311 );
    or g24690 ( n16904 , n13301 , n5528 );
    not g24691 ( n14010 , n14335 );
    not g24692 ( n27993 , n17968 );
    or g24693 ( n6120 , n13187 , n24450 );
    xnor g24694 ( n17660 , n2020 , n12116 );
    not g24695 ( n24539 , n12390 );
    nor g24696 ( n16582 , n27453 , n18518 );
    and g24697 ( n16530 , n29800 , n1572 );
    nor g24698 ( n30495 , n7983 , n11044 );
    xnor g24699 ( n12194 , n19894 , n18469 );
    xor g24700 ( n20577 , n20047 , n16052 );
    not g24701 ( n9200 , n24844 );
    or g24702 ( n30770 , n14860 , n3610 );
    and g24703 ( n8917 , n14098 , n28448 );
    not g24704 ( n2958 , n21584 );
    not g24705 ( n9053 , n30525 );
    not g24706 ( n22019 , n23232 );
    nor g24707 ( n10051 , n17918 , n7459 );
    xor g24708 ( n28724 , n27867 , n29974 );
    not g24709 ( n20366 , n17718 );
    nor g24710 ( n27679 , n2883 , n20822 );
    and g24711 ( n11586 , n23190 , n24746 );
    not g24712 ( n24934 , n16848 );
    or g24713 ( n4295 , n23097 , n15999 );
    xnor g24714 ( n15723 , n17138 , n25883 );
    xnor g24715 ( n31360 , n5827 , n20155 );
    xnor g24716 ( n8477 , n18190 , n27370 );
    nor g24717 ( n9019 , n6676 , n5550 );
    nor g24718 ( n1612 , n25841 , n18478 );
    not g24719 ( n20493 , n3101 );
    not g24720 ( n10480 , n17809 );
    not g24721 ( n16906 , n12086 );
    nor g24722 ( n30918 , n29298 , n16468 );
    or g24723 ( n19709 , n23364 , n7693 );
    xnor g24724 ( n25797 , n20846 , n859 );
    not g24725 ( n5336 , n22581 );
    or g24726 ( n22090 , n22747 , n25326 );
    and g24727 ( n24996 , n22108 , n30101 );
    xnor g24728 ( n18334 , n29124 , n26576 );
    xnor g24729 ( n12794 , n18970 , n7293 );
    and g24730 ( n2145 , n28737 , n17611 );
    and g24731 ( n12099 , n5128 , n397 );
    and g24732 ( n3162 , n23399 , n24690 );
    not g24733 ( n22775 , n22077 );
    not g24734 ( n29121 , n26867 );
    xnor g24735 ( n30634 , n13807 , n14683 );
    and g24736 ( n25564 , n10005 , n23287 );
    not g24737 ( n3514 , n25228 );
    not g24738 ( n27575 , n2570 );
    xor g24739 ( n13971 , n12780 , n16494 );
    xnor g24740 ( n23403 , n27395 , n6736 );
    and g24741 ( n14885 , n25451 , n21500 );
    and g24742 ( n13828 , n15033 , n27035 );
    not g24743 ( n19681 , n5854 );
    nor g24744 ( n11662 , n26863 , n9321 );
    or g24745 ( n15058 , n9486 , n6882 );
    xnor g24746 ( n10048 , n10071 , n20825 );
    xnor g24747 ( n1966 , n6811 , n9336 );
    nor g24748 ( n29703 , n31108 , n3289 );
    xnor g24749 ( n7232 , n25497 , n3677 );
    nor g24750 ( n12485 , n27435 , n10792 );
    or g24751 ( n25588 , n10838 , n24641 );
    xnor g24752 ( n23144 , n17614 , n30799 );
    nor g24753 ( n5767 , n4836 , n31847 );
    or g24754 ( n22995 , n2645 , n21637 );
    and g24755 ( n29633 , n31457 , n12442 );
    not g24756 ( n2701 , n18551 );
    and g24757 ( n829 , n26361 , n31429 );
    xnor g24758 ( n747 , n6593 , n16584 );
    or g24759 ( n26093 , n3335 , n3818 );
    xnor g24760 ( n19658 , n20453 , n2963 );
    or g24761 ( n27867 , n5783 , n15230 );
    and g24762 ( n22739 , n31932 , n972 );
    xnor g24763 ( n10820 , n14445 , n4393 );
    or g24764 ( n7430 , n31926 , n21188 );
    not g24765 ( n1380 , n4577 );
    and g24766 ( n30869 , n767 , n25623 );
    xnor g24767 ( n18023 , n29377 , n18865 );
    nor g24768 ( n18875 , n15010 , n11060 );
    or g24769 ( n23687 , n17859 , n23604 );
    xnor g24770 ( n928 , n23841 , n24849 );
    xnor g24771 ( n69 , n22083 , n2567 );
    or g24772 ( n11986 , n27917 , n21553 );
    not g24773 ( n8545 , n13627 );
    or g24774 ( n31349 , n3628 , n20898 );
    and g24775 ( n21181 , n19557 , n28065 );
    and g24776 ( n11606 , n27584 , n28284 );
    not g24777 ( n3072 , n1685 );
    not g24778 ( n9971 , n29424 );
    nor g24779 ( n3634 , n31201 , n11181 );
    xnor g24780 ( n1112 , n16722 , n31493 );
    not g24781 ( n977 , n21568 );
    not g24782 ( n21084 , n28490 );
    or g24783 ( n26851 , n31163 , n26160 );
    not g24784 ( n23588 , n26158 );
    and g24785 ( n4382 , n9506 , n10787 );
    or g24786 ( n5234 , n25106 , n13534 );
    or g24787 ( n30330 , n2572 , n2214 );
    not g24788 ( n9834 , n13918 );
    nor g24789 ( n4496 , n757 , n18491 );
    or g24790 ( n16554 , n26584 , n16465 );
    and g24791 ( n22403 , n7909 , n6041 );
    not g24792 ( n9150 , n16615 );
    not g24793 ( n1028 , n7465 );
    or g24794 ( n23322 , n3319 , n26669 );
    xnor g24795 ( n23870 , n25655 , n11539 );
    or g24796 ( n2349 , n11360 , n30067 );
    not g24797 ( n24361 , n9518 );
    xnor g24798 ( n23796 , n15255 , n9548 );
    or g24799 ( n24960 , n4583 , n6136 );
    not g24800 ( n6511 , n3278 );
    not g24801 ( n7988 , n29093 );
    or g24802 ( n24469 , n17259 , n11528 );
    nor g24803 ( n4584 , n26082 , n23342 );
    not g24804 ( n7471 , n5854 );
    or g24805 ( n7451 , n22641 , n28271 );
    or g24806 ( n23763 , n27731 , n17104 );
    or g24807 ( n31480 , n3075 , n28279 );
    not g24808 ( n12433 , n9374 );
    or g24809 ( n12885 , n10317 , n13489 );
    not g24810 ( n6634 , n16909 );
    or g24811 ( n21255 , n23099 , n26449 );
    not g24812 ( n27172 , n25334 );
    not g24813 ( n17739 , n11360 );
    nor g24814 ( n24702 , n11581 , n31729 );
    and g24815 ( n3368 , n23874 , n1332 );
    not g24816 ( n7762 , n10845 );
    not g24817 ( n20795 , n10734 );
    xnor g24818 ( n30540 , n11391 , n11792 );
    or g24819 ( n11707 , n26854 , n26533 );
    xor g24820 ( n30262 , n14217 , n350 );
    and g24821 ( n23700 , n10228 , n561 );
    and g24822 ( n31354 , n14723 , n18068 );
    xnor g24823 ( n4480 , n19818 , n24578 );
    xnor g24824 ( n8673 , n31070 , n11643 );
    not g24825 ( n8681 , n11706 );
    not g24826 ( n3584 , n3218 );
    nor g24827 ( n22250 , n3034 , n1783 );
    nor g24828 ( n18120 , n6839 , n15491 );
    not g24829 ( n14937 , n12182 );
    or g24830 ( n5718 , n19507 , n25110 );
    or g24831 ( n24075 , n10914 , n19804 );
    or g24832 ( n19984 , n27552 , n2515 );
    and g24833 ( n23573 , n22542 , n26189 );
    and g24834 ( n24366 , n8857 , n13978 );
    or g24835 ( n26192 , n2518 , n625 );
    xnor g24836 ( n10551 , n9897 , n9155 );
    not g24837 ( n17797 , n24537 );
    xnor g24838 ( n19976 , n14125 , n19361 );
    or g24839 ( n20624 , n14039 , n2704 );
    not g24840 ( n16362 , n3297 );
    xnor g24841 ( n27777 , n27848 , n24056 );
    xor g24842 ( n29566 , n29496 , n29159 );
    xnor g24843 ( n22089 , n4862 , n23469 );
    not g24844 ( n14679 , n213 );
    not g24845 ( n9904 , n24736 );
    or g24846 ( n29358 , n25014 , n13844 );
    xnor g24847 ( n30788 , n31932 , n19043 );
    not g24848 ( n25809 , n8449 );
    not g24849 ( n10773 , n29143 );
    or g24850 ( n28582 , n4924 , n29794 );
    and g24851 ( n18089 , n12482 , n4158 );
    not g24852 ( n7028 , n14035 );
    xnor g24853 ( n27278 , n2256 , n31696 );
    and g24854 ( n14701 , n12046 , n5464 );
    or g24855 ( n29612 , n30446 , n17728 );
    xnor g24856 ( n14978 , n861 , n4516 );
    not g24857 ( n12078 , n11755 );
    nor g24858 ( n9786 , n6300 , n820 );
    nor g24859 ( n29956 , n29726 , n6464 );
    xnor g24860 ( n3618 , n25277 , n10852 );
    not g24861 ( n4223 , n7594 );
    not g24862 ( n15612 , n18696 );
    or g24863 ( n728 , n31961 , n9923 );
    xnor g24864 ( n24598 , n10784 , n22140 );
    not g24865 ( n30793 , n4711 );
    and g24866 ( n28924 , n10500 , n16681 );
    nor g24867 ( n30385 , n29447 , n10897 );
    or g24868 ( n17384 , n27004 , n24669 );
    nor g24869 ( n7639 , n7821 , n1343 );
    or g24870 ( n30039 , n20584 , n13156 );
    or g24871 ( n14139 , n10295 , n1504 );
    not g24872 ( n20678 , n7731 );
    and g24873 ( n19395 , n6752 , n258 );
    not g24874 ( n8897 , n17019 );
    or g24875 ( n31645 , n13494 , n9443 );
    not g24876 ( n18525 , n31076 );
    not g24877 ( n5159 , n6659 );
    not g24878 ( n30471 , n4350 );
    not g24879 ( n11324 , n14069 );
    nor g24880 ( n15504 , n25089 , n29039 );
    or g24881 ( n4921 , n11075 , n21619 );
    not g24882 ( n19624 , n21465 );
    xnor g24883 ( n2824 , n14857 , n24513 );
    or g24884 ( n13537 , n10391 , n29516 );
    xnor g24885 ( n13092 , n24078 , n4235 );
    nor g24886 ( n10144 , n18558 , n9441 );
    or g24887 ( n3507 , n7412 , n27041 );
    not g24888 ( n27673 , n6923 );
    not g24889 ( n30037 , n3934 );
    nor g24890 ( n24605 , n7046 , n28245 );
    not g24891 ( n853 , n1524 );
    or g24892 ( n25876 , n4360 , n2507 );
    or g24893 ( n22513 , n20350 , n1294 );
    and g24894 ( n9963 , n23574 , n17319 );
    not g24895 ( n18543 , n469 );
    not g24896 ( n3611 , n26665 );
    or g24897 ( n10834 , n21422 , n31138 );
    and g24898 ( n8157 , n23138 , n24590 );
    or g24899 ( n22540 , n2040 , n22506 );
    not g24900 ( n26501 , n15692 );
    xnor g24901 ( n11206 , n3082 , n14714 );
    and g24902 ( n11830 , n31398 , n20737 );
    not g24903 ( n10147 , n8948 );
    xnor g24904 ( n1663 , n14589 , n29984 );
    nor g24905 ( n31577 , n10439 , n7896 );
    xnor g24906 ( n18586 , n829 , n31641 );
    and g24907 ( n30283 , n9917 , n3017 );
    xnor g24908 ( n17213 , n15378 , n15422 );
    xnor g24909 ( n23035 , n27017 , n1186 );
    or g24910 ( n28477 , n16193 , n15857 );
    xnor g24911 ( n23151 , n20374 , n508 );
    and g24912 ( n28393 , n21243 , n8713 );
    or g24913 ( n27400 , n27756 , n1171 );
    xor g24914 ( n5805 , n20144 , n26510 );
    xnor g24915 ( n20315 , n10592 , n17957 );
    and g24916 ( n18105 , n12702 , n28012 );
    not g24917 ( n15215 , n25882 );
    or g24918 ( n31597 , n31986 , n29319 );
    or g24919 ( n23918 , n14905 , n22834 );
    and g24920 ( n12501 , n8522 , n19864 );
    not g24921 ( n4421 , n23058 );
    xnor g24922 ( n27493 , n6905 , n14004 );
    buf g24923 ( n13939 , n25953 );
    nor g24924 ( n26775 , n31549 , n7799 );
    xnor g24925 ( n5066 , n8895 , n402 );
    not g24926 ( n18265 , n2998 );
    not g24927 ( n26710 , n31975 );
    xnor g24928 ( n6725 , n18854 , n345 );
    or g24929 ( n26497 , n27885 , n19113 );
    not g24930 ( n24201 , n21782 );
    xnor g24931 ( n25177 , n13505 , n31414 );
    or g24932 ( n8925 , n9134 , n12375 );
    xnor g24933 ( n3365 , n19172 , n8137 );
    or g24934 ( n25328 , n18130 , n2529 );
    or g24935 ( n29385 , n30529 , n27091 );
    xnor g24936 ( n15262 , n19158 , n29453 );
    xnor g24937 ( n20724 , n8544 , n25179 );
    not g24938 ( n27667 , n21708 );
    and g24939 ( n12176 , n14651 , n26457 );
    not g24940 ( n9269 , n3744 );
    or g24941 ( n6624 , n24056 , n29669 );
    and g24942 ( n27261 , n15837 , n31777 );
    xnor g24943 ( n18984 , n20072 , n32012 );
    nor g24944 ( n26911 , n28333 , n25409 );
    xnor g24945 ( n42 , n24299 , n3822 );
    not g24946 ( n10356 , n2359 );
    and g24947 ( n28142 , n6970 , n31727 );
    xor g24948 ( n7658 , n8807 , n29357 );
    and g24949 ( n5551 , n9914 , n6910 );
    not g24950 ( n31895 , n9693 );
    or g24951 ( n16297 , n8309 , n13564 );
    not g24952 ( n10862 , n2429 );
    or g24953 ( n20491 , n28634 , n21676 );
    and g24954 ( n26874 , n3496 , n14758 );
    not g24955 ( n13855 , n26424 );
    xnor g24956 ( n7854 , n23425 , n779 );
    not g24957 ( n13200 , n11321 );
    or g24958 ( n21763 , n26867 , n3412 );
    or g24959 ( n16027 , n27549 , n7933 );
    xnor g24960 ( n25624 , n14093 , n26768 );
    not g24961 ( n14993 , n31050 );
    not g24962 ( n26 , n4807 );
    or g24963 ( n10003 , n13822 , n28930 );
    nor g24964 ( n9863 , n31394 , n25392 );
    xnor g24965 ( n5457 , n19570 , n18645 );
    or g24966 ( n19148 , n9821 , n28460 );
    xnor g24967 ( n11500 , n1252 , n10794 );
    buf g24968 ( n19315 , n10774 );
    xnor g24969 ( n27497 , n7425 , n5069 );
    or g24970 ( n24972 , n23893 , n7205 );
    xnor g24971 ( n8093 , n24792 , n5022 );
    xnor g24972 ( n20050 , n748 , n6412 );
    or g24973 ( n27411 , n20770 , n1769 );
    not g24974 ( n13894 , n11366 );
    nor g24975 ( n4341 , n31727 , n21134 );
    xnor g24976 ( n13815 , n12865 , n19885 );
    xnor g24977 ( n16532 , n25226 , n26790 );
    xnor g24978 ( n13966 , n1720 , n21185 );
    xnor g24979 ( n20769 , n31867 , n4843 );
    or g24980 ( n30787 , n1195 , n27965 );
    or g24981 ( n20571 , n29216 , n11443 );
    xnor g24982 ( n24761 , n22300 , n10981 );
    or g24983 ( n9522 , n13724 , n14558 );
    or g24984 ( n336 , n17767 , n29778 );
    not g24985 ( n25851 , n10327 );
    and g24986 ( n12631 , n21296 , n12907 );
    not g24987 ( n15292 , n22994 );
    or g24988 ( n19060 , n4856 , n30886 );
    or g24989 ( n28827 , n573 , n21497 );
    and g24990 ( n6478 , n8237 , n1496 );
    or g24991 ( n18858 , n30627 , n12671 );
    not g24992 ( n16733 , n27933 );
    not g24993 ( n13138 , n10349 );
    xnor g24994 ( n14928 , n9463 , n29939 );
    xnor g24995 ( n6244 , n6371 , n23577 );
    xnor g24996 ( n26609 , n15562 , n24839 );
    nor g24997 ( n3286 , n22233 , n11674 );
    nor g24998 ( n16315 , n18391 , n6597 );
    xnor g24999 ( n28422 , n1081 , n20562 );
    or g25000 ( n18200 , n714 , n28088 );
    and g25001 ( n26364 , n16690 , n30514 );
    not g25002 ( n7775 , n4505 );
    not g25003 ( n14831 , n19617 );
    or g25004 ( n24133 , n8585 , n3141 );
    not g25005 ( n26728 , n6311 );
    and g25006 ( n12742 , n19297 , n11380 );
    not g25007 ( n2806 , n8969 );
    or g25008 ( n15743 , n18532 , n4638 );
    nor g25009 ( n603 , n1869 , n11976 );
    and g25010 ( n11628 , n18064 , n21990 );
    not g25011 ( n23125 , n8773 );
    xnor g25012 ( n1465 , n22255 , n3558 );
    not g25013 ( n31331 , n11900 );
    xnor g25014 ( n843 , n5022 , n19221 );
    nor g25015 ( n9023 , n26264 , n17380 );
    and g25016 ( n6432 , n26834 , n28350 );
    or g25017 ( n21045 , n25269 , n22687 );
    nor g25018 ( n10803 , n2924 , n17977 );
    or g25019 ( n11330 , n21708 , n19107 );
    nor g25020 ( n16731 , n20374 , n23433 );
    not g25021 ( n17322 , n5638 );
    and g25022 ( n10482 , n948 , n2386 );
    and g25023 ( n24523 , n26145 , n14594 );
    and g25024 ( n7429 , n6920 , n22651 );
    or g25025 ( n31598 , n20794 , n12345 );
    nor g25026 ( n9430 , n14544 , n3235 );
    xnor g25027 ( n26190 , n17693 , n22230 );
    not g25028 ( n27891 , n2825 );
    xnor g25029 ( n28537 , n14165 , n19424 );
    not g25030 ( n22119 , n30294 );
    not g25031 ( n23910 , n1476 );
    and g25032 ( n28480 , n23972 , n6341 );
    nor g25033 ( n27913 , n24152 , n20028 );
    or g25034 ( n23250 , n12696 , n23433 );
    xnor g25035 ( n30260 , n24791 , n27230 );
    or g25036 ( n11481 , n12122 , n16085 );
    xnor g25037 ( n26335 , n27209 , n9390 );
    or g25038 ( n13777 , n24185 , n3064 );
    or g25039 ( n22515 , n31338 , n12437 );
    nor g25040 ( n22360 , n16061 , n14206 );
    and g25041 ( n22213 , n21705 , n20710 );
    nor g25042 ( n17849 , n18761 , n21574 );
    and g25043 ( n3330 , n29687 , n21486 );
    xnor g25044 ( n27248 , n8001 , n11651 );
    not g25045 ( n25394 , n16152 );
    xnor g25046 ( n25930 , n26482 , n17039 );
    not g25047 ( n1299 , n22710 );
    and g25048 ( n25062 , n25752 , n176 );
    and g25049 ( n13421 , n1893 , n17279 );
    or g25050 ( n370 , n1333 , n14027 );
    and g25051 ( n25109 , n25301 , n7089 );
    not g25052 ( n13381 , n1692 );
    xnor g25053 ( n18148 , n18742 , n25416 );
    xnor g25054 ( n3905 , n20493 , n27113 );
    xnor g25055 ( n10956 , n11442 , n31069 );
    not g25056 ( n26327 , n11036 );
    not g25057 ( n15519 , n31386 );
    or g25058 ( n7906 , n13242 , n16914 );
    or g25059 ( n5107 , n32028 , n28002 );
    or g25060 ( n11844 , n5626 , n13907 );
    nor g25061 ( n22161 , n1728 , n19563 );
    and g25062 ( n16936 , n8913 , n20266 );
    nor g25063 ( n26177 , n22734 , n19474 );
    not g25064 ( n28091 , n19274 );
    not g25065 ( n12379 , n27064 );
    xnor g25066 ( n10996 , n15277 , n25630 );
    or g25067 ( n24493 , n11404 , n30869 );
    nor g25068 ( n19398 , n16299 , n906 );
    xnor g25069 ( n3722 , n3589 , n21700 );
    xnor g25070 ( n13737 , n16684 , n19425 );
    xnor g25071 ( n28606 , n4389 , n11131 );
    xnor g25072 ( n31637 , n10186 , n27888 );
    xnor g25073 ( n23832 , n11503 , n1231 );
    not g25074 ( n2570 , n17519 );
    xnor g25075 ( n20057 , n16666 , n9835 );
    and g25076 ( n7734 , n12560 , n30159 );
    and g25077 ( n2630 , n18100 , n31935 );
    and g25078 ( n7893 , n15515 , n29657 );
    or g25079 ( n29346 , n294 , n11951 );
    not g25080 ( n18869 , n26186 );
    not g25081 ( n9262 , n7180 );
    not g25082 ( n5237 , n11999 );
    nor g25083 ( n5620 , n17711 , n28034 );
    xnor g25084 ( n18432 , n28635 , n19211 );
    not g25085 ( n12086 , n23982 );
    or g25086 ( n22965 , n17579 , n30611 );
    and g25087 ( n28435 , n24538 , n5971 );
    not g25088 ( n1878 , n27334 );
    or g25089 ( n25117 , n15234 , n13290 );
    nor g25090 ( n28662 , n21272 , n12041 );
    or g25091 ( n10830 , n2093 , n25907 );
    not g25092 ( n10154 , n32010 );
    or g25093 ( n22990 , n26488 , n4146 );
    and g25094 ( n4191 , n8325 , n9748 );
    and g25095 ( n30507 , n9309 , n9076 );
    nor g25096 ( n23584 , n18234 , n16001 );
    and g25097 ( n30851 , n20037 , n5987 );
    and g25098 ( n11538 , n7066 , n18178 );
    xnor g25099 ( n5007 , n20849 , n3576 );
    and g25100 ( n29586 , n18366 , n20121 );
    not g25101 ( n25444 , n30389 );
    not g25102 ( n6780 , n20782 );
    xnor g25103 ( n1879 , n10037 , n26990 );
    not g25104 ( n21132 , n22454 );
    not g25105 ( n20660 , n8411 );
    xnor g25106 ( n22332 , n1938 , n10872 );
    or g25107 ( n30922 , n9969 , n4884 );
    and g25108 ( n13587 , n23442 , n304 );
    xnor g25109 ( n29359 , n6057 , n17920 );
    or g25110 ( n3211 , n7377 , n30639 );
    or g25111 ( n17702 , n20335 , n29714 );
    not g25112 ( n15981 , n22490 );
    not g25113 ( n17588 , n6199 );
    xnor g25114 ( n15043 , n10805 , n12857 );
    or g25115 ( n5164 , n20615 , n5115 );
    xnor g25116 ( n1467 , n2437 , n13711 );
    nor g25117 ( n14521 , n23040 , n29090 );
    not g25118 ( n5301 , n15132 );
    xnor g25119 ( n2047 , n7434 , n3076 );
    or g25120 ( n1162 , n11302 , n5143 );
    not g25121 ( n6063 , n23666 );
    and g25122 ( n29096 , n27300 , n16499 );
    not g25123 ( n1820 , n17620 );
    xnor g25124 ( n5385 , n27864 , n26068 );
    nor g25125 ( n14776 , n11691 , n15120 );
    not g25126 ( n28494 , n9912 );
    nor g25127 ( n11753 , n7033 , n7608 );
    or g25128 ( n15347 , n22314 , n21018 );
    or g25129 ( n12615 , n8426 , n1794 );
    xnor g25130 ( n22603 , n18099 , n48 );
    nor g25131 ( n29680 , n14913 , n12591 );
    not g25132 ( n22135 , n3500 );
    xor g25133 ( n3934 , n9658 , n29388 );
    not g25134 ( n19484 , n6111 );
    and g25135 ( n7956 , n14744 , n13974 );
    or g25136 ( n18892 , n19907 , n31520 );
    not g25137 ( n64 , n23218 );
    and g25138 ( n10277 , n28631 , n17061 );
    xnor g25139 ( n27996 , n25737 , n21402 );
    nor g25140 ( n31227 , n5752 , n8878 );
    not g25141 ( n10731 , n16414 );
    xnor g25142 ( n30276 , n31828 , n17370 );
    and g25143 ( n29877 , n12421 , n10567 );
    and g25144 ( n9750 , n14904 , n2463 );
    or g25145 ( n26672 , n20045 , n135 );
    nor g25146 ( n10711 , n6603 , n5305 );
    nor g25147 ( n18238 , n4526 , n18830 );
    and g25148 ( n16257 , n18673 , n14371 );
    not g25149 ( n10778 , n1212 );
    not g25150 ( n24164 , n20552 );
    or g25151 ( n14487 , n17194 , n31764 );
    and g25152 ( n23877 , n10830 , n22017 );
    not g25153 ( n12119 , n3531 );
    nor g25154 ( n14199 , n18394 , n16873 );
    or g25155 ( n13055 , n20008 , n8887 );
    not g25156 ( n11932 , n23614 );
    not g25157 ( n12711 , n15275 );
    not g25158 ( n29506 , n2454 );
    or g25159 ( n9125 , n5346 , n17121 );
    not g25160 ( n22718 , n14114 );
    and g25161 ( n18696 , n11806 , n18141 );
    not g25162 ( n17998 , n3473 );
    and g25163 ( n23385 , n15777 , n23210 );
    not g25164 ( n19777 , n13684 );
    xnor g25165 ( n25953 , n22506 , n24734 );
    nor g25166 ( n8981 , n25520 , n8291 );
    not g25167 ( n15887 , n12980 );
    not g25168 ( n29392 , n25636 );
    not g25169 ( n13552 , n4571 );
    xnor g25170 ( n5232 , n7612 , n22757 );
    or g25171 ( n31329 , n12754 , n14432 );
    xnor g25172 ( n18 , n26221 , n20278 );
    not g25173 ( n14646 , n14410 );
    not g25174 ( n14298 , n16655 );
    not g25175 ( n2657 , n28992 );
    not g25176 ( n14082 , n7604 );
    and g25177 ( n20938 , n29767 , n27870 );
    and g25178 ( n29516 , n19536 , n13766 );
    and g25179 ( n27475 , n1751 , n12514 );
    or g25180 ( n26166 , n25362 , n15273 );
    xnor g25181 ( n418 , n18078 , n23597 );
    not g25182 ( n23984 , n3272 );
    not g25183 ( n17515 , n2024 );
    not g25184 ( n27227 , n30562 );
    xnor g25185 ( n1865 , n6228 , n11996 );
    and g25186 ( n507 , n23841 , n24692 );
    not g25187 ( n3890 , n6318 );
    and g25188 ( n19975 , n18522 , n6013 );
    not g25189 ( n5473 , n10637 );
    nor g25190 ( n27385 , n31414 , n736 );
    or g25191 ( n5976 , n1195 , n22031 );
    not g25192 ( n1588 , n5037 );
    not g25193 ( n7580 , n7029 );
    or g25194 ( n20301 , n6394 , n7050 );
    nor g25195 ( n20784 , n10393 , n28258 );
    xnor g25196 ( n31287 , n30859 , n12449 );
    nor g25197 ( n3675 , n29351 , n1690 );
    not g25198 ( n19083 , n19959 );
    or g25199 ( n27593 , n4492 , n699 );
    not g25200 ( n1695 , n5103 );
    or g25201 ( n26946 , n1939 , n29013 );
    or g25202 ( n25080 , n28141 , n11491 );
    not g25203 ( n31592 , n6620 );
    not g25204 ( n13285 , n7775 );
    nor g25205 ( n9890 , n27000 , n17724 );
    and g25206 ( n6608 , n27128 , n31262 );
    and g25207 ( n32005 , n3325 , n7247 );
    nor g25208 ( n6945 , n29764 , n29604 );
    or g25209 ( n24432 , n2948 , n15079 );
    xnor g25210 ( n1818 , n14720 , n22574 );
    and g25211 ( n27788 , n18321 , n2935 );
    nor g25212 ( n16199 , n22316 , n25653 );
    nor g25213 ( n11697 , n27244 , n22707 );
    not g25214 ( n12066 , n3907 );
    not g25215 ( n24204 , n19883 );
    not g25216 ( n21633 , n10699 );
    or g25217 ( n11678 , n15883 , n6173 );
    nor g25218 ( n29556 , n2432 , n17820 );
    xnor g25219 ( n24500 , n8647 , n24118 );
    or g25220 ( n2157 , n22427 , n1548 );
    xnor g25221 ( n14743 , n761 , n6722 );
    not g25222 ( n1585 , n5255 );
    or g25223 ( n6303 , n9712 , n23080 );
    not g25224 ( n16476 , n15619 );
    xnor g25225 ( n5122 , n10034 , n30505 );
    or g25226 ( n4893 , n2630 , n6868 );
    not g25227 ( n3383 , n13527 );
    or g25228 ( n23849 , n31409 , n14284 );
    and g25229 ( n7317 , n27696 , n1367 );
    nor g25230 ( n21491 , n11488 , n9745 );
    xnor g25231 ( n4663 , n21802 , n19873 );
    nor g25232 ( n2436 , n19125 , n19084 );
    or g25233 ( n10280 , n2758 , n18732 );
    or g25234 ( n31441 , n26842 , n17280 );
    and g25235 ( n16940 , n4803 , n20038 );
    xnor g25236 ( n5564 , n5569 , n20677 );
    or g25237 ( n9355 , n24166 , n31388 );
    xnor g25238 ( n31693 , n5808 , n25797 );
    and g25239 ( n30783 , n18858 , n25568 );
    not g25240 ( n20402 , n4316 );
    and g25241 ( n10396 , n23645 , n17186 );
    and g25242 ( n24836 , n12538 , n273 );
    not g25243 ( n12170 , n3281 );
    nor g25244 ( n13628 , n14521 , n17431 );
    xnor g25245 ( n21688 , n11977 , n13090 );
    not g25246 ( n14844 , n1699 );
    nor g25247 ( n7810 , n97 , n10451 );
    xnor g25248 ( n9673 , n29732 , n4032 );
    or g25249 ( n2921 , n16538 , n25681 );
    and g25250 ( n25986 , n17389 , n3814 );
    and g25251 ( n11805 , n969 , n29881 );
    xnor g25252 ( n8324 , n29224 , n29615 );
    or g25253 ( n28312 , n1990 , n9858 );
    or g25254 ( n27003 , n14715 , n9890 );
    not g25255 ( n10017 , n3288 );
    not g25256 ( n27732 , n29721 );
    and g25257 ( n25979 , n20460 , n28591 );
    not g25258 ( n11043 , n29143 );
    xnor g25259 ( n29148 , n17965 , n29655 );
    and g25260 ( n15528 , n15001 , n27156 );
    and g25261 ( n2121 , n30475 , n2152 );
    or g25262 ( n31944 , n26118 , n22397 );
    xnor g25263 ( n19620 , n17022 , n16450 );
    xnor g25264 ( n10004 , n20886 , n12729 );
    nor g25265 ( n6914 , n5237 , n12790 );
    xnor g25266 ( n18867 , n15019 , n10122 );
    not g25267 ( n15097 , n21029 );
    xnor g25268 ( n19823 , n12850 , n21980 );
    or g25269 ( n19015 , n2482 , n15264 );
    xnor g25270 ( n17462 , n10050 , n7026 );
    nor g25271 ( n29473 , n7784 , n10666 );
    or g25272 ( n12748 , n24939 , n7028 );
    not g25273 ( n16011 , n19474 );
    not g25274 ( n10044 , n21089 );
    not g25275 ( n22930 , n26873 );
    not g25276 ( n23119 , n16132 );
    xnor g25277 ( n21459 , n9228 , n22451 );
    and g25278 ( n19216 , n17698 , n24886 );
    or g25279 ( n21848 , n26718 , n24655 );
    xnor g25280 ( n28804 , n28928 , n15572 );
    not g25281 ( n10473 , n5600 );
    xnor g25282 ( n27672 , n30417 , n3580 );
    xnor g25283 ( n29024 , n30411 , n26082 );
    or g25284 ( n17419 , n23986 , n21818 );
    or g25285 ( n5692 , n30620 , n18824 );
    or g25286 ( n11410 , n31406 , n761 );
    or g25287 ( n2892 , n4859 , n5564 );
    or g25288 ( n8997 , n13549 , n24826 );
    or g25289 ( n16173 , n20400 , n17111 );
    or g25290 ( n1605 , n17869 , n24499 );
    xnor g25291 ( n7674 , n19572 , n3108 );
    not g25292 ( n14704 , n21122 );
    nor g25293 ( n10503 , n5388 , n10327 );
    not g25294 ( n29642 , n1830 );
    not g25295 ( n12474 , n12607 );
    xnor g25296 ( n1012 , n17431 , n28155 );
    not g25297 ( n25201 , n13170 );
    nor g25298 ( n22199 , n22522 , n11868 );
    and g25299 ( n1998 , n8554 , n3474 );
    xnor g25300 ( n16701 , n14488 , n24961 );
    not g25301 ( n16871 , n11052 );
    and g25302 ( n2852 , n16021 , n26105 );
    not g25303 ( n952 , n31032 );
    and g25304 ( n27183 , n27535 , n5559 );
    not g25305 ( n12685 , n10120 );
    nor g25306 ( n16565 , n24569 , n27420 );
    and g25307 ( n7815 , n15766 , n7712 );
    and g25308 ( n1171 , n8615 , n728 );
    not g25309 ( n5563 , n1518 );
    xnor g25310 ( n22091 , n13370 , n25601 );
    not g25311 ( n19861 , n28794 );
    not g25312 ( n1535 , n4041 );
    or g25313 ( n27543 , n14420 , n21641 );
    or g25314 ( n6049 , n30340 , n5079 );
    xnor g25315 ( n10487 , n7973 , n11752 );
    xnor g25316 ( n4729 , n13791 , n7465 );
    and g25317 ( n1223 , n19766 , n6463 );
    nor g25318 ( n21100 , n14555 , n26032 );
    nor g25319 ( n18062 , n7564 , n21029 );
    xnor g25320 ( n29037 , n30171 , n7789 );
    not g25321 ( n15398 , n4542 );
    not g25322 ( n6165 , n13614 );
    xnor g25323 ( n27041 , n27697 , n12360 );
    or g25324 ( n22311 , n23755 , n28097 );
    nor g25325 ( n19121 , n25793 , n15122 );
    not g25326 ( n18751 , n13758 );
    xnor g25327 ( n18529 , n28266 , n18890 );
    and g25328 ( n26738 , n11122 , n31137 );
    not g25329 ( n31106 , n5022 );
    or g25330 ( n3294 , n25163 , n15117 );
    and g25331 ( n4137 , n29286 , n6606 );
    not g25332 ( n31905 , n10627 );
    or g25333 ( n1726 , n5359 , n25575 );
    and g25334 ( n25003 , n8599 , n24603 );
    not g25335 ( n24678 , n2323 );
    nor g25336 ( n1053 , n13957 , n606 );
    or g25337 ( n22183 , n10308 , n4879 );
    nor g25338 ( n12037 , n13020 , n31817 );
    and g25339 ( n12228 , n24646 , n17621 );
    and g25340 ( n19012 , n23952 , n6231 );
    or g25341 ( n9867 , n30632 , n12564 );
    or g25342 ( n27871 , n15887 , n28061 );
    or g25343 ( n18016 , n17283 , n22485 );
    or g25344 ( n3794 , n770 , n4752 );
    xnor g25345 ( n1422 , n21587 , n24748 );
    and g25346 ( n23602 , n29352 , n15707 );
    and g25347 ( n7819 , n26829 , n2500 );
    and g25348 ( n13905 , n23526 , n40 );
    xnor g25349 ( n31802 , n6495 , n31352 );
    xnor g25350 ( n5201 , n16159 , n31153 );
    not g25351 ( n25414 , n17057 );
    and g25352 ( n15419 , n1560 , n17188 );
    not g25353 ( n30555 , n24435 );
    or g25354 ( n19994 , n6652 , n2321 );
    not g25355 ( n21428 , n29315 );
    xnor g25356 ( n19949 , n16336 , n21510 );
    xnor g25357 ( n16670 , n13855 , n25212 );
    xnor g25358 ( n23275 , n4916 , n10120 );
    or g25359 ( n28352 , n3591 , n10105 );
    xnor g25360 ( n5727 , n22707 , n13849 );
    or g25361 ( n29884 , n9414 , n17037 );
    not g25362 ( n11980 , n30579 );
    not g25363 ( n26397 , n19198 );
    not g25364 ( n16202 , n6849 );
    nor g25365 ( n10030 , n5712 , n31821 );
    and g25366 ( n10523 , n29338 , n8074 );
    xnor g25367 ( n6880 , n7349 , n13417 );
    xnor g25368 ( n21873 , n6721 , n8862 );
    xnor g25369 ( n4673 , n17812 , n30343 );
    and g25370 ( n22614 , n29104 , n22980 );
    not g25371 ( n21687 , n24613 );
    xnor g25372 ( n11035 , n23609 , n12948 );
    buf g25373 ( n2200 , n459 );
    and g25374 ( n8495 , n1041 , n15352 );
    and g25375 ( n4289 , n31117 , n26770 );
    not g25376 ( n21871 , n28828 );
    xnor g25377 ( n3425 , n25247 , n15458 );
    not g25378 ( n6346 , n238 );
    or g25379 ( n2350 , n1962 , n27250 );
    or g25380 ( n24296 , n4582 , n20326 );
    not g25381 ( n13415 , n11763 );
    xnor g25382 ( n30929 , n9935 , n19217 );
    nor g25383 ( n20417 , n494 , n19067 );
    not g25384 ( n22025 , n1194 );
    or g25385 ( n9305 , n3641 , n27965 );
    or g25386 ( n27225 , n27505 , n28971 );
    and g25387 ( n17678 , n24357 , n21830 );
    xnor g25388 ( n10823 , n21242 , n10196 );
    not g25389 ( n21769 , n4305 );
    not g25390 ( n19571 , n11069 );
    not g25391 ( n10507 , n9596 );
    not g25392 ( n22169 , n24360 );
    nor g25393 ( n25804 , n7927 , n30991 );
    not g25394 ( n27929 , n11246 );
    and g25395 ( n4879 , n20542 , n94 );
    not g25396 ( n608 , n20803 );
    nor g25397 ( n23396 , n23669 , n22129 );
    and g25398 ( n8244 , n15039 , n30203 );
    or g25399 ( n23969 , n21094 , n13789 );
    not g25400 ( n29807 , n19233 );
    nor g25401 ( n14416 , n29663 , n2097 );
    xnor g25402 ( n16900 , n18169 , n17333 );
    or g25403 ( n1157 , n23176 , n30196 );
    or g25404 ( n23473 , n21993 , n17714 );
    or g25405 ( n25240 , n8470 , n30816 );
    or g25406 ( n4156 , n27900 , n16316 );
    not g25407 ( n21789 , n26996 );
    xnor g25408 ( n27960 , n11223 , n9209 );
    xnor g25409 ( n16003 , n8186 , n22466 );
    nor g25410 ( n9389 , n8978 , n22935 );
    or g25411 ( n3188 , n17784 , n7385 );
    not g25412 ( n6009 , n14090 );
    xnor g25413 ( n5141 , n29917 , n17857 );
    not g25414 ( n27000 , n12605 );
    not g25415 ( n17985 , n4779 );
    and g25416 ( n15308 , n17908 , n9521 );
    and g25417 ( n29899 , n640 , n14389 );
    not g25418 ( n14812 , n31309 );
    not g25419 ( n16633 , n7707 );
    or g25420 ( n8016 , n5150 , n1889 );
    and g25421 ( n12614 , n9319 , n9320 );
    or g25422 ( n9309 , n2776 , n7329 );
    and g25423 ( n13190 , n30619 , n5107 );
    not g25424 ( n15866 , n21284 );
    xnor g25425 ( n7518 , n30530 , n20632 );
    or g25426 ( n28456 , n13976 , n12690 );
    xor g25427 ( n19196 , n4083 , n226 );
    not g25428 ( n19236 , n10151 );
    xnor g25429 ( n29831 , n31855 , n13318 );
    and g25430 ( n6814 , n4666 , n845 );
    not g25431 ( n8252 , n30160 );
    not g25432 ( n22204 , n17491 );
    buf g25433 ( n29879 , n8475 );
    or g25434 ( n25345 , n18326 , n9110 );
    not g25435 ( n9162 , n3793 );
    or g25436 ( n11757 , n17035 , n25168 );
    and g25437 ( n10988 , n25221 , n25494 );
    xnor g25438 ( n14110 , n29537 , n9697 );
    not g25439 ( n9849 , n18744 );
    xnor g25440 ( n26518 , n18071 , n20504 );
    or g25441 ( n13133 , n18825 , n17130 );
    nor g25442 ( n31958 , n28758 , n10188 );
    xnor g25443 ( n8087 , n7461 , n27449 );
    not g25444 ( n4704 , n12772 );
    xnor g25445 ( n4445 , n2249 , n18880 );
    not g25446 ( n2221 , n28035 );
    xnor g25447 ( n10763 , n24052 , n22681 );
    and g25448 ( n25127 , n3034 , n26512 );
    nor g25449 ( n8996 , n31970 , n5654 );
    xnor g25450 ( n4568 , n11399 , n13598 );
    or g25451 ( n6805 , n15469 , n30051 );
    and g25452 ( n24655 , n8793 , n31207 );
    and g25453 ( n5490 , n9758 , n21312 );
    not g25454 ( n3709 , n31325 );
    and g25455 ( n1046 , n22202 , n11155 );
    and g25456 ( n10916 , n22273 , n25561 );
    or g25457 ( n29488 , n21230 , n8059 );
    not g25458 ( n26511 , n28270 );
    xnor g25459 ( n6192 , n23184 , n12207 );
    xnor g25460 ( n4887 , n12690 , n19333 );
    xnor g25461 ( n8869 , n15134 , n4379 );
    xnor g25462 ( n25369 , n3368 , n24500 );
    not g25463 ( n25358 , n3426 );
    xor g25464 ( n19188 , n23713 , n25793 );
    not g25465 ( n24153 , n4742 );
    or g25466 ( n15653 , n5121 , n13446 );
    not g25467 ( n11298 , n28920 );
    not g25468 ( n6277 , n24522 );
    buf g25469 ( n11028 , n22411 );
    xnor g25470 ( n21569 , n24659 , n15780 );
    not g25471 ( n23999 , n25763 );
    or g25472 ( n29730 , n31580 , n9462 );
    and g25473 ( n21915 , n28190 , n23233 );
    not g25474 ( n29870 , n30187 );
    and g25475 ( n13483 , n20513 , n13557 );
    or g25476 ( n21618 , n6044 , n27573 );
    not g25477 ( n2085 , n826 );
    or g25478 ( n1912 , n572 , n18501 );
    and g25479 ( n18109 , n21214 , n18965 );
    not g25480 ( n15365 , n9136 );
    nor g25481 ( n17877 , n21300 , n13818 );
    not g25482 ( n31393 , n5697 );
    xnor g25483 ( n9680 , n3654 , n28859 );
    and g25484 ( n8065 , n15757 , n19341 );
    nor g25485 ( n6297 , n8808 , n12055 );
    or g25486 ( n10000 , n30918 , n31886 );
    nor g25487 ( n17741 , n10740 , n4665 );
    or g25488 ( n10766 , n26234 , n15942 );
    or g25489 ( n17792 , n26095 , n30055 );
    or g25490 ( n9253 , n11325 , n10876 );
    xnor g25491 ( n8118 , n26750 , n18762 );
    not g25492 ( n4789 , n7209 );
    or g25493 ( n19674 , n26125 , n26475 );
    xnor g25494 ( n27030 , n8440 , n5501 );
    and g25495 ( n821 , n21215 , n24976 );
    nor g25496 ( n4098 , n8321 , n29134 );
    xnor g25497 ( n3293 , n13268 , n20486 );
    not g25498 ( n28164 , n18867 );
    not g25499 ( n30433 , n5396 );
    or g25500 ( n27100 , n19030 , n24864 );
    or g25501 ( n10998 , n20514 , n30707 );
    nor g25502 ( n16620 , n22107 , n15928 );
    xnor g25503 ( n23379 , n26967 , n28938 );
    xnor g25504 ( n24206 , n29668 , n24415 );
    nor g25505 ( n30791 , n22174 , n2177 );
    not g25506 ( n9596 , n13075 );
    xnor g25507 ( n19869 , n10158 , n30458 );
    xnor g25508 ( n7987 , n24729 , n23448 );
    or g25509 ( n12447 , n20857 , n10593 );
    not g25510 ( n8896 , n29686 );
    not g25511 ( n24420 , n13338 );
    or g25512 ( n5910 , n3940 , n25375 );
    nor g25513 ( n31409 , n9520 , n17746 );
    not g25514 ( n20436 , n12727 );
    not g25515 ( n15301 , n624 );
    not g25516 ( n25196 , n14507 );
    and g25517 ( n6953 , n20581 , n12611 );
    xnor g25518 ( n21442 , n18172 , n4296 );
    xnor g25519 ( n5459 , n23737 , n18690 );
    not g25520 ( n24254 , n20713 );
    or g25521 ( n890 , n1953 , n1107 );
    or g25522 ( n13246 , n28417 , n1204 );
    not g25523 ( n25454 , n17628 );
    or g25524 ( n20719 , n3731 , n7068 );
    nor g25525 ( n17332 , n28709 , n7424 );
    xnor g25526 ( n30971 , n987 , n1301 );
    not g25527 ( n16421 , n21301 );
    xnor g25528 ( n2536 , n5558 , n6196 );
    not g25529 ( n20554 , n26783 );
    nor g25530 ( n27527 , n1177 , n28136 );
    not g25531 ( n30366 , n17430 );
    xnor g25532 ( n28460 , n29906 , n11218 );
    xor g25533 ( n27275 , n12053 , n24377 );
    or g25534 ( n30101 , n1194 , n18311 );
    nor g25535 ( n28648 , n23852 , n28562 );
    or g25536 ( n11099 , n12788 , n17190 );
    and g25537 ( n18136 , n24096 , n16502 );
    not g25538 ( n11123 , n25543 );
    xnor g25539 ( n20125 , n25541 , n12242 );
    and g25540 ( n5491 , n28849 , n23459 );
    and g25541 ( n16983 , n17297 , n9379 );
    and g25542 ( n5702 , n29211 , n29277 );
    xnor g25543 ( n3651 , n28015 , n2649 );
    xnor g25544 ( n7168 , n16277 , n6256 );
    not g25545 ( n10155 , n29114 );
    nor g25546 ( n26539 , n8364 , n19852 );
    xnor g25547 ( n19208 , n19997 , n22228 );
    xnor g25548 ( n21832 , n30686 , n17652 );
    and g25549 ( n30981 , n3181 , n20422 );
    and g25550 ( n25823 , n18256 , n6413 );
    not g25551 ( n25130 , n1692 );
    or g25552 ( n26803 , n16741 , n25887 );
    xnor g25553 ( n13177 , n6167 , n16216 );
    xnor g25554 ( n1531 , n11213 , n16287 );
    or g25555 ( n8614 , n30805 , n24724 );
    not g25556 ( n7118 , n9402 );
    xnor g25557 ( n23453 , n21857 , n16210 );
    xor g25558 ( n10853 , n28110 , n10670 );
    or g25559 ( n22629 , n27778 , n31130 );
    not g25560 ( n15062 , n19967 );
    and g25561 ( n19677 , n19225 , n20592 );
    xnor g25562 ( n21615 , n11365 , n8214 );
    xnor g25563 ( n7583 , n6175 , n17390 );
    xnor g25564 ( n11770 , n11488 , n6554 );
    xor g25565 ( n23611 , n24497 , n6224 );
    and g25566 ( n31537 , n19582 , n14846 );
    xnor g25567 ( n1849 , n12021 , n6848 );
    or g25568 ( n2465 , n24132 , n7514 );
    nor g25569 ( n31384 , n11866 , n31783 );
    and g25570 ( n18942 , n8339 , n15596 );
    not g25571 ( n3462 , n16672 );
    not g25572 ( n1920 , n27253 );
    xnor g25573 ( n24494 , n9730 , n27322 );
    or g25574 ( n1620 , n23218 , n30706 );
    xnor g25575 ( n26345 , n8258 , n3786 );
    or g25576 ( n7550 , n22172 , n17602 );
    not g25577 ( n1418 , n12448 );
    and g25578 ( n25584 , n30823 , n24343 );
    not g25579 ( n13081 , n1555 );
    or g25580 ( n4279 , n12030 , n17558 );
    xnor g25581 ( n18288 , n12281 , n20088 );
    xnor g25582 ( n4829 , n21466 , n17995 );
    xnor g25583 ( n4510 , n21562 , n17895 );
    and g25584 ( n27256 , n20298 , n26772 );
    not g25585 ( n14042 , n29961 );
    and g25586 ( n31024 , n9214 , n9405 );
    xnor g25587 ( n5963 , n12040 , n13498 );
    not g25588 ( n15794 , n9121 );
    xnor g25589 ( n29238 , n4731 , n9752 );
    not g25590 ( n8971 , n31303 );
    or g25591 ( n15316 , n10949 , n1853 );
    not g25592 ( n29290 , n423 );
    and g25593 ( n2757 , n13508 , n20815 );
    xnor g25594 ( n25491 , n21481 , n31266 );
    xnor g25595 ( n24803 , n7057 , n31190 );
    not g25596 ( n15517 , n27650 );
    not g25597 ( n7908 , n3804 );
    not g25598 ( n21941 , n17910 );
    or g25599 ( n31300 , n1421 , n21987 );
    xnor g25600 ( n14968 , n30706 , n13859 );
    or g25601 ( n21802 , n19081 , n29928 );
    not g25602 ( n10137 , n1415 );
    not g25603 ( n30950 , n2727 );
    or g25604 ( n25073 , n5531 , n12045 );
    or g25605 ( n12442 , n24455 , n21708 );
    and g25606 ( n1682 , n16547 , n23228 );
    not g25607 ( n29403 , n10636 );
    and g25608 ( n12109 , n21446 , n17177 );
    not g25609 ( n18559 , n25397 );
    xor g25610 ( n23962 , n19241 , n4179 );
    not g25611 ( n30293 , n29171 );
    or g25612 ( n16636 , n10469 , n2747 );
    not g25613 ( n30795 , n14184 );
    xnor g25614 ( n27448 , n19096 , n31143 );
    xnor g25615 ( n31907 , n23216 , n12660 );
    not g25616 ( n3012 , n23236 );
    or g25617 ( n3865 , n5856 , n24869 );
    not g25618 ( n20327 , n828 );
    and g25619 ( n10344 , n31463 , n13284 );
    and g25620 ( n18971 , n21149 , n15212 );
    xnor g25621 ( n9406 , n10214 , n20019 );
    or g25622 ( n16665 , n3570 , n12004 );
    xnor g25623 ( n31173 , n4541 , n19625 );
    or g25624 ( n10425 , n12300 , n18747 );
    not g25625 ( n31754 , n31104 );
    xnor g25626 ( n29075 , n14508 , n5831 );
    not g25627 ( n26823 , n3837 );
    or g25628 ( n24123 , n14884 , n27834 );
    not g25629 ( n1582 , n3719 );
    xnor g25630 ( n28514 , n21528 , n11012 );
    and g25631 ( n8850 , n13469 , n12120 );
    nor g25632 ( n23846 , n23179 , n24972 );
    buf g25633 ( n953 , n4459 );
    xnor g25634 ( n509 , n16203 , n23145 );
    not g25635 ( n1821 , n3996 );
    and g25636 ( n17214 , n8272 , n7085 );
    not g25637 ( n21741 , n23870 );
    or g25638 ( n6064 , n18953 , n19714 );
    and g25639 ( n76 , n13408 , n27551 );
    and g25640 ( n14465 , n5705 , n3807 );
    not g25641 ( n8945 , n19939 );
    xnor g25642 ( n4631 , n23529 , n11928 );
    not g25643 ( n8603 , n792 );
    or g25644 ( n12000 , n32008 , n20427 );
    xnor g25645 ( n26267 , n14020 , n20805 );
    and g25646 ( n2525 , n26496 , n16729 );
    xnor g25647 ( n4108 , n8139 , n27002 );
    or g25648 ( n6844 , n25231 , n12269 );
    and g25649 ( n30286 , n4744 , n18667 );
    not g25650 ( n11990 , n30057 );
    xnor g25651 ( n20410 , n27588 , n25877 );
    and g25652 ( n11108 , n25902 , n14690 );
    or g25653 ( n22782 , n17197 , n13693 );
    not g25654 ( n28885 , n121 );
    xor g25655 ( n2529 , n7673 , n13835 );
    xnor g25656 ( n23499 , n1860 , n11360 );
    not g25657 ( n4079 , n18979 );
    xnor g25658 ( n26585 , n15020 , n5299 );
    and g25659 ( n9897 , n30718 , n9630 );
    and g25660 ( n26490 , n16339 , n16410 );
    not g25661 ( n13590 , n18816 );
    xnor g25662 ( n11281 , n27934 , n12262 );
    not g25663 ( n4835 , n25350 );
    or g25664 ( n11509 , n6476 , n9365 );
    nor g25665 ( n1128 , n6145 , n5294 );
    nor g25666 ( n25149 , n19956 , n138 );
    or g25667 ( n30778 , n2226 , n6308 );
    xnor g25668 ( n20826 , n10126 , n16765 );
    not g25669 ( n11717 , n22339 );
    or g25670 ( n23625 , n9299 , n25973 );
    or g25671 ( n6017 , n31964 , n20947 );
    not g25672 ( n16078 , n5362 );
    and g25673 ( n22566 , n19520 , n24749 );
    xnor g25674 ( n25200 , n1922 , n30897 );
    xnor g25675 ( n18959 , n12990 , n22248 );
    xnor g25676 ( n16398 , n30730 , n3336 );
    xnor g25677 ( n28069 , n1336 , n9781 );
    nor g25678 ( n22018 , n22973 , n13477 );
    not g25679 ( n24948 , n20569 );
    and g25680 ( n15216 , n2592 , n15382 );
    nor g25681 ( n28274 , n12920 , n19675 );
    not g25682 ( n23449 , n31966 );
    and g25683 ( n18084 , n30454 , n13000 );
    not g25684 ( n20226 , n12582 );
    or g25685 ( n26917 , n19428 , n15523 );
    nor g25686 ( n11700 , n16103 , n16373 );
    xnor g25687 ( n28212 , n14760 , n12617 );
    and g25688 ( n744 , n16553 , n17594 );
    or g25689 ( n14818 , n4274 , n18068 );
    not g25690 ( n15573 , n8875 );
    and g25691 ( n19686 , n26985 , n20166 );
    not g25692 ( n2220 , n8910 );
    xnor g25693 ( n2861 , n24525 , n11643 );
    or g25694 ( n4436 , n10957 , n6573 );
    or g25695 ( n26416 , n13737 , n29871 );
    nor g25696 ( n30155 , n11692 , n6757 );
    xnor g25697 ( n28671 , n22569 , n14792 );
    not g25698 ( n25435 , n30976 );
    or g25699 ( n2468 , n14222 , n21226 );
    xnor g25700 ( n969 , n31175 , n4651 );
    not g25701 ( n24230 , n14492 );
    not g25702 ( n11763 , n9259 );
    not g25703 ( n23967 , n31218 );
    and g25704 ( n23237 , n20908 , n25313 );
    not g25705 ( n3111 , n4997 );
    and g25706 ( n22285 , n20136 , n20375 );
    and g25707 ( n26903 , n4679 , n935 );
    nor g25708 ( n22818 , n18551 , n12777 );
    not g25709 ( n18465 , n12812 );
    not g25710 ( n7355 , n30002 );
    not g25711 ( n26386 , n18462 );
    not g25712 ( n11694 , n11453 );
    xnor g25713 ( n3066 , n6078 , n20427 );
    not g25714 ( n16782 , n16534 );
    nor g25715 ( n31919 , n13170 , n3505 );
    nor g25716 ( n661 , n4599 , n704 );
    xnor g25717 ( n11273 , n25760 , n13454 );
    not g25718 ( n2490 , n7932 );
    nor g25719 ( n23188 , n28774 , n12203 );
    or g25720 ( n3705 , n1608 , n10387 );
    and g25721 ( n23664 , n13832 , n2099 );
    nor g25722 ( n20329 , n6871 , n18895 );
    not g25723 ( n9211 , n18730 );
    xnor g25724 ( n4275 , n1341 , n17640 );
    not g25725 ( n27555 , n10845 );
    not g25726 ( n20303 , n13869 );
    or g25727 ( n9332 , n25161 , n30488 );
    or g25728 ( n4825 , n28205 , n9960 );
    not g25729 ( n27706 , n23608 );
    xnor g25730 ( n21780 , n23196 , n12509 );
    xnor g25731 ( n3746 , n4778 , n18170 );
    nor g25732 ( n21478 , n594 , n12961 );
    not g25733 ( n21436 , n25680 );
    not g25734 ( n6738 , n27960 );
    nor g25735 ( n2915 , n31651 , n2437 );
    or g25736 ( n1715 , n30579 , n5503 );
    not g25737 ( n14669 , n8081 );
    xnor g25738 ( n1784 , n5746 , n12803 );
    not g25739 ( n26365 , n12732 );
    not g25740 ( n30935 , n27770 );
    xnor g25741 ( n4926 , n16050 , n4661 );
    not g25742 ( n26137 , n24153 );
    nor g25743 ( n15296 , n10071 , n25793 );
    and g25744 ( n12192 , n9035 , n23289 );
    and g25745 ( n4261 , n6303 , n26847 );
    and g25746 ( n194 , n19978 , n21839 );
    or g25747 ( n12651 , n16764 , n120 );
    and g25748 ( n11469 , n19227 , n10601 );
    not g25749 ( n6585 , n15619 );
    not g25750 ( n435 , n8903 );
    not g25751 ( n22031 , n18362 );
    not g25752 ( n7851 , n22594 );
    xnor g25753 ( n22807 , n14382 , n14408 );
    xnor g25754 ( n11760 , n19528 , n20358 );
    not g25755 ( n10366 , n25271 );
    not g25756 ( n25674 , n25117 );
    and g25757 ( n18472 , n12842 , n23250 );
    and g25758 ( n18154 , n307 , n5584 );
    not g25759 ( n10423 , n22549 );
    nor g25760 ( n19088 , n11658 , n12602 );
    or g25761 ( n23623 , n5966 , n15456 );
    xnor g25762 ( n22141 , n29209 , n16670 );
    not g25763 ( n16975 , n24250 );
    or g25764 ( n11828 , n25092 , n4777 );
    nor g25765 ( n20672 , n17363 , n30982 );
    not g25766 ( n23523 , n9059 );
    xnor g25767 ( n300 , n19314 , n4257 );
    xnor g25768 ( n18788 , n2123 , n13472 );
    not g25769 ( n25687 , n31185 );
    nor g25770 ( n6806 , n22169 , n13029 );
    xnor g25771 ( n8625 , n11746 , n14504 );
    xnor g25772 ( n18718 , n8005 , n30411 );
    xor g25773 ( n26185 , n28679 , n7014 );
    not g25774 ( n17217 , n29290 );
    nor g25775 ( n23251 , n28983 , n4246 );
    xnor g25776 ( n11405 , n3810 , n17417 );
    not g25777 ( n16478 , n14134 );
    not g25778 ( n28341 , n2798 );
    not g25779 ( n5882 , n4830 );
    xnor g25780 ( n3815 , n12959 , n30813 );
    nor g25781 ( n31145 , n11500 , n2126 );
    not g25782 ( n16076 , n25137 );
    xor g25783 ( n26494 , n22115 , n20664 );
    not g25784 ( n11220 , n1516 );
    and g25785 ( n24888 , n12197 , n19180 );
    not g25786 ( n930 , n30273 );
    nor g25787 ( n751 , n25318 , n1241 );
    xnor g25788 ( n5496 , n15420 , n29593 );
    or g25789 ( n4857 , n7102 , n6580 );
    xnor g25790 ( n1073 , n29562 , n2335 );
    or g25791 ( n18738 , n3688 , n8283 );
    xnor g25792 ( n28300 , n7463 , n24286 );
    xnor g25793 ( n15944 , n17391 , n7896 );
    and g25794 ( n12902 , n16979 , n23855 );
    xnor g25795 ( n12126 , n29486 , n27541 );
    or g25796 ( n15643 , n30458 , n20536 );
    or g25797 ( n25834 , n1626 , n11096 );
    not g25798 ( n5132 , n6789 );
    or g25799 ( n3650 , n20284 , n21352 );
    xnor g25800 ( n18857 , n13231 , n7272 );
    or g25801 ( n26442 , n29370 , n3316 );
    nor g25802 ( n22683 , n25210 , n25915 );
    and g25803 ( n30446 , n22545 , n31516 );
    or g25804 ( n11078 , n2712 , n20233 );
    not g25805 ( n340 , n19679 );
    or g25806 ( n16696 , n4522 , n30730 );
    not g25807 ( n2889 , n29201 );
    and g25808 ( n22565 , n19996 , n14322 );
    or g25809 ( n20119 , n5280 , n21435 );
    or g25810 ( n26189 , n25334 , n4054 );
    xnor g25811 ( n20330 , n30238 , n11643 );
    not g25812 ( n25871 , n16858 );
    nor g25813 ( n26171 , n20510 , n27227 );
    xnor g25814 ( n27694 , n20916 , n20038 );
    xnor g25815 ( n7539 , n16466 , n18947 );
    xnor g25816 ( n15988 , n2302 , n29797 );
    or g25817 ( n7215 , n11953 , n17848 );
    xnor g25818 ( n13521 , n31520 , n2370 );
    not g25819 ( n8516 , n17497 );
    not g25820 ( n1482 , n12061 );
    not g25821 ( n15899 , n14924 );
    nor g25822 ( n26089 , n24522 , n21982 );
    xnor g25823 ( n27434 , n26636 , n24056 );
    or g25824 ( n4444 , n12520 , n11150 );
    or g25825 ( n2419 , n8315 , n22285 );
    not g25826 ( n9625 , n21931 );
    nor g25827 ( n6682 , n8308 , n2679 );
    and g25828 ( n22767 , n23847 , n27423 );
    and g25829 ( n17077 , n15345 , n20026 );
    xnor g25830 ( n6462 , n28573 , n11025 );
    or g25831 ( n22955 , n4097 , n25109 );
    xnor g25832 ( n10734 , n24231 , n9400 );
    or g25833 ( n27938 , n7675 , n10066 );
    nor g25834 ( n24124 , n15999 , n7414 );
    and g25835 ( n31984 , n29917 , n8248 );
    and g25836 ( n18323 , n25910 , n23363 );
    or g25837 ( n21939 , n28177 , n19687 );
    xnor g25838 ( n16191 , n25608 , n29116 );
    xnor g25839 ( n12264 , n26862 , n28435 );
    and g25840 ( n16969 , n18796 , n17485 );
    not g25841 ( n1704 , n12988 );
    not g25842 ( n14513 , n17499 );
    not g25843 ( n30112 , n2483 );
    or g25844 ( n4782 , n24415 , n20708 );
    or g25845 ( n11337 , n11587 , n1049 );
    nor g25846 ( n15761 , n14711 , n6871 );
    not g25847 ( n23624 , n12776 );
    and g25848 ( n10078 , n20852 , n20370 );
    not g25849 ( n2070 , n29418 );
    xnor g25850 ( n11461 , n3808 , n23423 );
    not g25851 ( n2599 , n24003 );
    or g25852 ( n29722 , n97 , n11880 );
    not g25853 ( n3848 , n23856 );
    and g25854 ( n9167 , n22569 , n14792 );
    nor g25855 ( n25833 , n11890 , n2389 );
    and g25856 ( n7326 , n14622 , n13340 );
    buf g25857 ( n1366 , n15991 );
    not g25858 ( n6406 , n14063 );
    not g25859 ( n18972 , n27550 );
    nor g25860 ( n20347 , n9831 , n7745 );
    or g25861 ( n16832 , n19692 , n6472 );
    xnor g25862 ( n13594 , n144 , n17107 );
    and g25863 ( n19682 , n12789 , n15978 );
    or g25864 ( n1835 , n29377 , n7170 );
    xnor g25865 ( n4783 , n25455 , n12766 );
    or g25866 ( n14500 , n7703 , n30496 );
    and g25867 ( n10230 , n23412 , n9466 );
    not g25868 ( n10454 , n7491 );
    not g25869 ( n15724 , n18060 );
    xnor g25870 ( n1593 , n30500 , n14273 );
    not g25871 ( n12759 , n16524 );
    or g25872 ( n12413 , n9239 , n9362 );
    xnor g25873 ( n28931 , n21280 , n8196 );
    xnor g25874 ( n7736 , n21998 , n674 );
    or g25875 ( n23797 , n2601 , n28573 );
    or g25876 ( n15383 , n27447 , n6589 );
    or g25877 ( n31872 , n14679 , n24766 );
    not g25878 ( n18074 , n28712 );
    not g25879 ( n17363 , n6446 );
    or g25880 ( n21211 , n4415 , n16648 );
    xnor g25881 ( n20382 , n2905 , n21191 );
    xnor g25882 ( n25680 , n5667 , n31212 );
    and g25883 ( n21523 , n6361 , n22652 );
    not g25884 ( n12641 , n5833 );
    and g25885 ( n19948 , n21975 , n27076 );
    and g25886 ( n25307 , n11460 , n17277 );
    or g25887 ( n9972 , n21516 , n16819 );
    xnor g25888 ( n305 , n445 , n2883 );
    not g25889 ( n20920 , n28633 );
    xnor g25890 ( n21332 , n20121 , n21407 );
    xnor g25891 ( n22773 , n12927 , n17776 );
    not g25892 ( n14713 , n31544 );
    or g25893 ( n5644 , n25680 , n5272 );
    or g25894 ( n23381 , n31082 , n13486 );
    xnor g25895 ( n1495 , n8578 , n7701 );
    or g25896 ( n23227 , n14824 , n4186 );
    xnor g25897 ( n1144 , n8155 , n29320 );
    and g25898 ( n2364 , n11335 , n29509 );
    or g25899 ( n7885 , n3214 , n4592 );
    or g25900 ( n16745 , n9370 , n3955 );
    xnor g25901 ( n8836 , n4546 , n3063 );
    nor g25902 ( n31280 , n26823 , n20252 );
    not g25903 ( n4644 , n25679 );
    or g25904 ( n29597 , n12399 , n9135 );
    buf g25905 ( n6696 , n29261 );
    xnor g25906 ( n22277 , n9028 , n24601 );
    xnor g25907 ( n15325 , n17704 , n22916 );
    or g25908 ( n6991 , n24837 , n23115 );
    and g25909 ( n8518 , n19647 , n24907 );
    or g25910 ( n16337 , n14072 , n10999 );
    or g25911 ( n18175 , n4386 , n31243 );
    and g25912 ( n25241 , n7561 , n17522 );
    or g25913 ( n23989 , n18653 , n16155 );
    or g25914 ( n30395 , n12515 , n31046 );
    or g25915 ( n5035 , n11315 , n8179 );
    not g25916 ( n1891 , n13494 );
    buf g25917 ( n5834 , n25978 );
    xnor g25918 ( n12076 , n24512 , n16799 );
    xnor g25919 ( n12136 , n23056 , n18955 );
    xnor g25920 ( n12500 , n22634 , n7090 );
    not g25921 ( n30190 , n19488 );
    not g25922 ( n17766 , n15391 );
    not g25923 ( n15636 , n6676 );
    and g25924 ( n31242 , n9489 , n11009 );
    or g25925 ( n27934 , n30818 , n10472 );
    or g25926 ( n31554 , n10864 , n11697 );
    or g25927 ( n28732 , n29132 , n25403 );
    and g25928 ( n7454 , n29868 , n5195 );
    xnor g25929 ( n27939 , n26456 , n12514 );
    or g25930 ( n18480 , n13323 , n18592 );
    xnor g25931 ( n6168 , n28042 , n29086 );
    or g25932 ( n14186 , n27074 , n24205 );
    not g25933 ( n5746 , n2574 );
    or g25934 ( n16634 , n5153 , n1324 );
    xnor g25935 ( n8270 , n10212 , n616 );
    xor g25936 ( n12856 , n28686 , n9636 );
    or g25937 ( n3324 , n10389 , n10097 );
    or g25938 ( n8205 , n31475 , n1998 );
    not g25939 ( n5912 , n16368 );
    and g25940 ( n7912 , n29244 , n3764 );
    or g25941 ( n23654 , n26504 , n9114 );
    and g25942 ( n19209 , n17996 , n12177 );
    xnor g25943 ( n21700 , n27594 , n27529 );
    xnor g25944 ( n27705 , n23843 , n31878 );
    not g25945 ( n24128 , n7216 );
    xnor g25946 ( n21866 , n21711 , n6957 );
    xnor g25947 ( n5897 , n24440 , n7707 );
    xnor g25948 ( n21748 , n19145 , n4131 );
    not g25949 ( n850 , n16414 );
    xnor g25950 ( n4845 , n8713 , n11065 );
    or g25951 ( n20091 , n6309 , n31935 );
    or g25952 ( n31504 , n15307 , n23063 );
    xnor g25953 ( n16278 , n11611 , n6696 );
    xnor g25954 ( n1897 , n20614 , n16981 );
    not g25955 ( n386 , n28632 );
    xnor g25956 ( n13689 , n15758 , n17843 );
    and g25957 ( n23300 , n28061 , n1178 );
    not g25958 ( n25791 , n4257 );
    or g25959 ( n22518 , n13131 , n22189 );
    and g25960 ( n17815 , n23774 , n16255 );
    not g25961 ( n28198 , n18130 );
    xnor g25962 ( n4917 , n9871 , n28494 );
    and g25963 ( n15169 , n1835 , n27102 );
    or g25964 ( n24344 , n793 , n1339 );
    nor g25965 ( n31613 , n30374 , n21158 );
    not g25966 ( n22857 , n810 );
    or g25967 ( n17188 , n25774 , n20360 );
    or g25968 ( n21776 , n31060 , n22233 );
    not g25969 ( n30476 , n18706 );
    or g25970 ( n22964 , n28682 , n16050 );
    and g25971 ( n26535 , n646 , n6250 );
    not g25972 ( n28314 , n7314 );
    or g25973 ( n5821 , n25215 , n16530 );
    or g25974 ( n28641 , n2618 , n16299 );
    or g25975 ( n9188 , n31016 , n10212 );
    and g25976 ( n9346 , n4564 , n22258 );
    xnor g25977 ( n14004 , n14080 , n21765 );
    or g25978 ( n20355 , n29238 , n8731 );
    and g25979 ( n9858 , n19015 , n30354 );
    xnor g25980 ( n18035 , n29633 , n16491 );
    or g25981 ( n24159 , n30129 , n27771 );
    and g25982 ( n28548 , n10769 , n238 );
    xnor g25983 ( n11366 , n19547 , n25361 );
    xnor g25984 ( n3578 , n15219 , n1997 );
    not g25985 ( n28627 , n17080 );
    not g25986 ( n14681 , n11327 );
    and g25987 ( n16396 , n24862 , n25073 );
    or g25988 ( n21095 , n23206 , n19744 );
    or g25989 ( n27297 , n28313 , n31451 );
    not g25990 ( n15808 , n23673 );
    or g25991 ( n27840 , n14117 , n4692 );
    xnor g25992 ( n6150 , n1328 , n24601 );
    or g25993 ( n9564 , n30697 , n17253 );
    xnor g25994 ( n2245 , n31282 , n26517 );
    not g25995 ( n29475 , n3449 );
    not g25996 ( n5809 , n10569 );
    not g25997 ( n12411 , n9625 );
    not g25998 ( n7576 , n20881 );
    not g25999 ( n18562 , n7313 );
    and g26000 ( n15670 , n2534 , n11483 );
    xnor g26001 ( n10056 , n25588 , n7422 );
    xnor g26002 ( n25137 , n22822 , n15933 );
    not g26003 ( n5153 , n442 );
    and g26004 ( n14223 , n9415 , n5021 );
    or g26005 ( n6876 , n27219 , n5309 );
    not g26006 ( n31033 , n26616 );
    xnor g26007 ( n21420 , n10749 , n1592 );
    and g26008 ( n22168 , n457 , n30749 );
    nor g26009 ( n30315 , n1217 , n3082 );
    nor g26010 ( n26095 , n9971 , n2882 );
    xnor g26011 ( n5880 , n2247 , n21006 );
    or g26012 ( n20429 , n17201 , n2123 );
    nor g26013 ( n8660 , n25699 , n17051 );
    not g26014 ( n22255 , n3359 );
    and g26015 ( n14226 , n4437 , n24176 );
    and g26016 ( n7597 , n28014 , n30824 );
    not g26017 ( n27352 , n4124 );
    or g26018 ( n19723 , n16421 , n787 );
    and g26019 ( n13595 , n25522 , n27509 );
    or g26020 ( n3020 , n21376 , n28602 );
    or g26021 ( n21481 , n7827 , n75 );
    or g26022 ( n8751 , n9939 , n11711 );
    or g26023 ( n24106 , n20799 , n11947 );
    not g26024 ( n6873 , n12392 );
    or g26025 ( n22992 , n20720 , n12472 );
    and g26026 ( n3528 , n22950 , n4481 );
    not g26027 ( n28068 , n14055 );
    or g26028 ( n28064 , n9777 , n26637 );
    not g26029 ( n27055 , n259 );
    nor g26030 ( n13727 , n22549 , n17499 );
    xnor g26031 ( n8028 , n14555 , n16200 );
    not g26032 ( n18922 , n20262 );
    xnor g26033 ( n21385 , n16219 , n30347 );
    xnor g26034 ( n2994 , n26609 , n21186 );
    not g26035 ( n4779 , n17357 );
    or g26036 ( n755 , n13401 , n21318 );
    and g26037 ( n3856 , n3222 , n25435 );
    and g26038 ( n9402 , n21988 , n15844 );
    xnor g26039 ( n5641 , n4803 , n26165 );
    nor g26040 ( n10006 , n12668 , n18506 );
    and g26041 ( n3610 , n8651 , n3671 );
    and g26042 ( n10720 , n25138 , n16143 );
    xnor g26043 ( n26159 , n8808 , n12055 );
    or g26044 ( n23009 , n29495 , n27424 );
    not g26045 ( n20015 , n22254 );
    or g26046 ( n29181 , n16664 , n24017 );
    not g26047 ( n14269 , n28756 );
    or g26048 ( n19774 , n128 , n29977 );
    not g26049 ( n26934 , n30306 );
    or g26050 ( n28229 , n15504 , n13862 );
    xnor g26051 ( n12390 , n4284 , n6096 );
    xnor g26052 ( n2400 , n16796 , n1630 );
    or g26053 ( n1070 , n5316 , n10733 );
    and g26054 ( n12019 , n11784 , n4099 );
    and g26055 ( n28363 , n26264 , n29567 );
    or g26056 ( n7233 , n31029 , n6530 );
    and g26057 ( n26664 , n13923 , n14967 );
    not g26058 ( n3430 , n5991 );
    xnor g26059 ( n22521 , n4717 , n30470 );
    or g26060 ( n26370 , n30287 , n22210 );
    nor g26061 ( n2309 , n7425 , n5069 );
    or g26062 ( n3739 , n13825 , n5176 );
    xnor g26063 ( n25172 , n13409 , n13102 );
    xnor g26064 ( n25673 , n26146 , n6680 );
    and g26065 ( n8488 , n27671 , n1513 );
    xnor g26066 ( n16511 , n23242 , n29576 );
    xnor g26067 ( n694 , n19211 , n7707 );
    and g26068 ( n12873 , n17392 , n8884 );
    xnor g26069 ( n10127 , n14052 , n12804 );
    or g26070 ( n23812 , n12516 , n7617 );
    not g26071 ( n11972 , n2617 );
    not g26072 ( n7526 , n26467 );
    not g26073 ( n7765 , n2444 );
    not g26074 ( n2017 , n8507 );
    or g26075 ( n1149 , n2222 , n27481 );
    and g26076 ( n30295 , n25152 , n13838 );
    nor g26077 ( n651 , n31812 , n23292 );
    xnor g26078 ( n13249 , n699 , n19731 );
    and g26079 ( n20288 , n18615 , n15287 );
    and g26080 ( n19494 , n21194 , n5296 );
    nor g26081 ( n21536 , n4161 , n22814 );
    not g26082 ( n777 , n6938 );
    xnor g26083 ( n12570 , n12308 , n22841 );
    or g26084 ( n1374 , n18106 , n26250 );
    xnor g26085 ( n5650 , n21379 , n8434 );
    and g26086 ( n9701 , n24779 , n7850 );
    not g26087 ( n10321 , n19159 );
    xnor g26088 ( n6883 , n877 , n3774 );
    xnor g26089 ( n20977 , n30022 , n12806 );
    xnor g26090 ( n19394 , n7271 , n5672 );
    xnor g26091 ( n28599 , n6528 , n22256 );
    xnor g26092 ( n4977 , n6527 , n31108 );
    not g26093 ( n3512 , n7682 );
    xnor g26094 ( n15030 , n19562 , n29572 );
    or g26095 ( n22492 , n20249 , n27928 );
    xnor g26096 ( n1713 , n26004 , n23342 );
    and g26097 ( n9432 , n22888 , n17397 );
    xnor g26098 ( n10388 , n31950 , n8593 );
    xnor g26099 ( n17023 , n18780 , n30245 );
    not g26100 ( n2993 , n22620 );
    xnor g26101 ( n13910 , n19175 , n8515 );
    xnor g26102 ( n29144 , n26191 , n10949 );
    and g26103 ( n29719 , n8383 , n23792 );
    nor g26104 ( n31163 , n16978 , n22022 );
    xnor g26105 ( n10768 , n21987 , n381 );
    or g26106 ( n30539 , n29635 , n7932 );
    nor g26107 ( n468 , n28686 , n4678 );
    or g26108 ( n31893 , n2904 , n26635 );
    xnor g26109 ( n14714 , n2150 , n11065 );
    xnor g26110 ( n1973 , n30843 , n12877 );
    not g26111 ( n9206 , n7417 );
    xnor g26112 ( n13925 , n19615 , n3614 );
    not g26113 ( n28652 , n18625 );
    not g26114 ( n27758 , n11035 );
    xnor g26115 ( n6833 , n27069 , n5924 );
    nor g26116 ( n2755 , n9642 , n25601 );
    or g26117 ( n15267 , n18262 , n25782 );
    xnor g26118 ( n23204 , n21838 , n12699 );
    nor g26119 ( n30128 , n995 , n23459 );
    and g26120 ( n7249 , n21900 , n27624 );
    xnor g26121 ( n28551 , n18631 , n1671 );
    nor g26122 ( n23534 , n1318 , n18605 );
    not g26123 ( n25403 , n561 );
    and g26124 ( n6540 , n4768 , n23943 );
    not g26125 ( n12130 , n25536 );
    or g26126 ( n23710 , n6148 , n3005 );
    nor g26127 ( n15644 , n13764 , n28179 );
    not g26128 ( n25818 , n22316 );
    not g26129 ( n2739 , n29520 );
    and g26130 ( n20553 , n16253 , n1838 );
    or g26131 ( n8146 , n6130 , n4454 );
    xnor g26132 ( n5625 , n1252 , n9826 );
    xnor g26133 ( n6862 , n23593 , n5533 );
    xnor g26134 ( n4209 , n5322 , n16978 );
    or g26135 ( n11806 , n29703 , n30780 );
    xnor g26136 ( n16755 , n18135 , n16799 );
    and g26137 ( n28204 , n27511 , n14106 );
    or g26138 ( n19277 , n601 , n26921 );
    xnor g26139 ( n19481 , n13046 , n16815 );
    not g26140 ( n25727 , n11694 );
    not g26141 ( n26654 , n10636 );
    xnor g26142 ( n21665 , n107 , n30458 );
    xnor g26143 ( n29470 , n15469 , n24716 );
    xnor g26144 ( n18392 , n17176 , n14477 );
    xnor g26145 ( n13886 , n20378 , n24588 );
    xnor g26146 ( n19421 , n28306 , n31918 );
    or g26147 ( n15368 , n13335 , n27514 );
    and g26148 ( n18554 , n12835 , n22034 );
    xnor g26149 ( n12888 , n9366 , n16579 );
    buf g26150 ( n7026 , n16858 );
    xnor g26151 ( n584 , n1039 , n10474 );
    xnor g26152 ( n11822 , n2430 , n16398 );
    or g26153 ( n28469 , n30272 , n22761 );
    xnor g26154 ( n24315 , n4844 , n27233 );
    xnor g26155 ( n21979 , n25271 , n15805 );
    not g26156 ( n27961 , n11178 );
    xnor g26157 ( n11506 , n12628 , n4924 );
    xor g26158 ( n10701 , n22395 , n17910 );
    xnor g26159 ( n19759 , n19015 , n24891 );
    xnor g26160 ( n6414 , n1517 , n23148 );
    and g26161 ( n17681 , n15477 , n30440 );
    or g26162 ( n15285 , n10857 , n3177 );
    nor g26163 ( n27717 , n7659 , n16709 );
    xnor g26164 ( n29846 , n28106 , n84 );
    not g26165 ( n26373 , n7046 );
    xnor g26166 ( n4555 , n27957 , n16833 );
    and g26167 ( n24155 , n13413 , n11065 );
    not g26168 ( n6015 , n14709 );
    or g26169 ( n17286 , n19977 , n23624 );
    not g26170 ( n31028 , n26368 );
    xnor g26171 ( n8057 , n20830 , n19206 );
    xnor g26172 ( n8536 , n18740 , n3494 );
    xnor g26173 ( n24540 , n25776 , n23195 );
    and g26174 ( n4676 , n1098 , n17051 );
    or g26175 ( n12208 , n3110 , n11924 );
    and g26176 ( n26663 , n20775 , n9892 );
    and g26177 ( n8665 , n10217 , n15184 );
    or g26178 ( n12218 , n15182 , n19948 );
    or g26179 ( n30802 , n19217 , n12198 );
    or g26180 ( n10761 , n16558 , n26073 );
    and g26181 ( n2942 , n14508 , n18210 );
    or g26182 ( n20370 , n31492 , n25290 );
    not g26183 ( n27532 , n15345 );
    not g26184 ( n31969 , n30706 );
    not g26185 ( n7391 , n31301 );
    nor g26186 ( n15137 , n18647 , n7787 );
    buf g26187 ( n21381 , n26943 );
    not g26188 ( n29499 , n25917 );
    not g26189 ( n25900 , n30505 );
    not g26190 ( n1707 , n25173 );
    not g26191 ( n20583 , n19615 );
    or g26192 ( n18811 , n12101 , n16612 );
    not g26193 ( n9485 , n2993 );
    and g26194 ( n18411 , n9147 , n28227 );
    xnor g26195 ( n18094 , n18391 , n9619 );
    not g26196 ( n24782 , n12511 );
    xnor g26197 ( n14683 , n18420 , n1045 );
    not g26198 ( n24397 , n110 );
    and g26199 ( n18815 , n20353 , n28841 );
    not g26200 ( n27550 , n3645 );
    or g26201 ( n21770 , n16411 , n25818 );
    or g26202 ( n4263 , n7210 , n17558 );
    and g26203 ( n26283 , n2363 , n18039 );
    and g26204 ( n1087 , n6351 , n27110 );
    xnor g26205 ( n4710 , n3787 , n18730 );
    not g26206 ( n14975 , n15162 );
    or g26207 ( n27923 , n30813 , n31563 );
    and g26208 ( n12852 , n18927 , n28477 );
    not g26209 ( n263 , n28210 );
    or g26210 ( n30110 , n17149 , n7576 );
    nor g26211 ( n10539 , n7593 , n1097 );
    and g26212 ( n430 , n18887 , n16912 );
    xnor g26213 ( n30656 , n3824 , n12425 );
    or g26214 ( n16258 , n31611 , n23039 );
    xnor g26215 ( n1687 , n17544 , n23905 );
    or g26216 ( n10128 , n16975 , n27474 );
    and g26217 ( n5663 , n8653 , n23531 );
    xnor g26218 ( n23502 , n23136 , n7902 );
    or g26219 ( n17938 , n27440 , n12976 );
    and g26220 ( n9426 , n28976 , n4409 );
    or g26221 ( n8697 , n11759 , n30494 );
    or g26222 ( n29619 , n21872 , n1622 );
    xnor g26223 ( n26914 , n1063 , n20168 );
    not g26224 ( n17310 , n13518 );
    xnor g26225 ( n22762 , n15682 , n12431 );
    or g26226 ( n23564 , n16758 , n4613 );
    nor g26227 ( n3042 , n27132 , n16302 );
    xnor g26228 ( n21624 , n7939 , n20561 );
    not g26229 ( n4577 , n14050 );
    xnor g26230 ( n8522 , n18426 , n14569 );
    or g26231 ( n17341 , n23159 , n11571 );
    xnor g26232 ( n14243 , n27217 , n23774 );
    xnor g26233 ( n29050 , n6121 , n6560 );
    or g26234 ( n22309 , n26607 , n10904 );
    xor g26235 ( n2723 , n7873 , n2262 );
    not g26236 ( n23340 , n24431 );
    not g26237 ( n1667 , n25247 );
    or g26238 ( n25667 , n10617 , n3245 );
    or g26239 ( n30001 , n15394 , n30097 );
    xnor g26240 ( n14049 , n11219 , n7093 );
    and g26241 ( n3589 , n10149 , n1342 );
    not g26242 ( n21374 , n19456 );
    or g26243 ( n363 , n22825 , n14395 );
    not g26244 ( n19717 , n11238 );
    and g26245 ( n13091 , n2505 , n31164 );
    nor g26246 ( n23971 , n20902 , n2294 );
    and g26247 ( n4129 , n447 , n18033 );
    xnor g26248 ( n21390 , n10761 , n17617 );
    and g26249 ( n30375 , n28382 , n22978 );
    and g26250 ( n950 , n19185 , n11361 );
    or g26251 ( n18937 , n10369 , n6400 );
    not g26252 ( n16174 , n11506 );
    or g26253 ( n8206 , n26036 , n25036 );
    nor g26254 ( n26112 , n23658 , n31719 );
    and g26255 ( n20634 , n18569 , n15551 );
    or g26256 ( n10517 , n16725 , n29560 );
    nor g26257 ( n23018 , n11060 , n26988 );
    not g26258 ( n13250 , n21709 );
    xnor g26259 ( n23311 , n18201 , n28387 );
    or g26260 ( n16463 , n1233 , n10462 );
    not g26261 ( n20209 , n22393 );
    not g26262 ( n4541 , n3676 );
    not g26263 ( n19292 , n7574 );
    not g26264 ( n27166 , n21646 );
    xnor g26265 ( n18373 , n17647 , n30514 );
    not g26266 ( n31369 , n1119 );
    or g26267 ( n14331 , n13328 , n5339 );
    nor g26268 ( n19612 , n20736 , n19871 );
    not g26269 ( n28689 , n2610 );
    nor g26270 ( n10566 , n26237 , n13184 );
    nor g26271 ( n4657 , n26052 , n13110 );
    and g26272 ( n30173 , n24826 , n13549 );
    not g26273 ( n26247 , n29132 );
    not g26274 ( n30895 , n24102 );
    not g26275 ( n21297 , n11360 );
    not g26276 ( n11598 , n31819 );
    xnor g26277 ( n30111 , n16323 , n20555 );
    not g26278 ( n15224 , n31954 );
    or g26279 ( n11544 , n757 , n14601 );
    not g26280 ( n26389 , n2018 );
    or g26281 ( n17553 , n1740 , n20033 );
    xnor g26282 ( n24895 , n19180 , n7881 );
    xnor g26283 ( n17242 , n3379 , n13583 );
    xnor g26284 ( n17207 , n9744 , n15010 );
    xnor g26285 ( n22121 , n11397 , n3019 );
    not g26286 ( n100 , n30964 );
    xnor g26287 ( n20291 , n8942 , n14116 );
    xnor g26288 ( n29524 , n29444 , n29974 );
    not g26289 ( n26290 , n11896 );
    xnor g26290 ( n24675 , n16519 , n4621 );
    xnor g26291 ( n24648 , n10564 , n15523 );
    not g26292 ( n9495 , n5020 );
    and g26293 ( n24091 , n21721 , n5605 );
    not g26294 ( n10002 , n15030 );
    xnor g26295 ( n21783 , n11026 , n26921 );
    not g26296 ( n24695 , n12772 );
    or g26297 ( n4633 , n19502 , n802 );
    and g26298 ( n29200 , n16221 , n9352 );
    xnor g26299 ( n8570 , n23006 , n8132 );
    xnor g26300 ( n17498 , n8904 , n15943 );
    or g26301 ( n21839 , n717 , n1699 );
    and g26302 ( n2557 , n12823 , n14440 );
    xor g26303 ( n18236 , n27963 , n24578 );
    xnor g26304 ( n17883 , n30870 , n23275 );
    not g26305 ( n29323 , n727 );
    not g26306 ( n10755 , n10643 );
    or g26307 ( n9979 , n2144 , n20047 );
    not g26308 ( n16461 , n4886 );
    or g26309 ( n3549 , n1262 , n7227 );
    not g26310 ( n20839 , n19747 );
    or g26311 ( n5591 , n11140 , n27438 );
    xnor g26312 ( n9322 , n12478 , n16019 );
    not g26313 ( n18264 , n24289 );
    not g26314 ( n3372 , n14557 );
    not g26315 ( n15056 , n27143 );
    xnor g26316 ( n3698 , n24367 , n18005 );
    or g26317 ( n30413 , n30034 , n11923 );
    not g26318 ( n9152 , n31864 );
    xnor g26319 ( n15791 , n30403 , n24651 );
    not g26320 ( n13431 , n24110 );
    not g26321 ( n13113 , n364 );
    nor g26322 ( n31053 , n22806 , n596 );
    and g26323 ( n30185 , n9146 , n11894 );
    and g26324 ( n23636 , n9631 , n26222 );
    or g26325 ( n23054 , n20978 , n14939 );
    or g26326 ( n12869 , n1809 , n9108 );
    xnor g26327 ( n31076 , n5513 , n16072 );
    xnor g26328 ( n2255 , n955 , n26008 );
    nor g26329 ( n5043 , n25610 , n25398 );
    and g26330 ( n22959 , n5335 , n19219 );
    or g26331 ( n10992 , n8416 , n9738 );
    nor g26332 ( n11210 , n2635 , n8103 );
    and g26333 ( n19816 , n23338 , n17266 );
    not g26334 ( n18611 , n12036 );
    or g26335 ( n3109 , n12232 , n12624 );
    not g26336 ( n16221 , n13433 );
    or g26337 ( n11480 , n22665 , n18360 );
    xnor g26338 ( n32012 , n17910 , n7655 );
    and g26339 ( n23973 , n18390 , n4677 );
    or g26340 ( n25853 , n25748 , n29712 );
    and g26341 ( n15247 , n13891 , n414 );
    xnor g26342 ( n12127 , n15903 , n30742 );
    or g26343 ( n22698 , n11290 , n26269 );
    and g26344 ( n18830 , n27869 , n15368 );
    or g26345 ( n29863 , n25077 , n8461 );
    not g26346 ( n17711 , n18617 );
    not g26347 ( n11561 , n5455 );
    not g26348 ( n11466 , n28562 );
    and g26349 ( n3087 , n26376 , n19218 );
    xnor g26350 ( n17665 , n20848 , n22244 );
    xnor g26351 ( n24610 , n8893 , n7017 );
    nor g26352 ( n4371 , n1 , n18524 );
    or g26353 ( n8203 , n17556 , n6730 );
    not g26354 ( n20588 , n5585 );
    or g26355 ( n14709 , n10213 , n5378 );
    or g26356 ( n26673 , n12574 , n14505 );
    not g26357 ( n27514 , n15291 );
    xor g26358 ( n17899 , n3364 , n9939 );
    not g26359 ( n22202 , n16281 );
    not g26360 ( n29407 , n11504 );
    xnor g26361 ( n23310 , n31261 , n18867 );
    or g26362 ( n6548 , n2565 , n7815 );
    xnor g26363 ( n4675 , n28224 , n922 );
    nor g26364 ( n6782 , n31894 , n25198 );
    not g26365 ( n14239 , n31790 );
    and g26366 ( n31943 , n29799 , n20300 );
    or g26367 ( n23746 , n14828 , n11324 );
    xnor g26368 ( n3252 , n27453 , n18518 );
    not g26369 ( n16292 , n2933 );
    or g26370 ( n16095 , n29346 , n23505 );
    xnor g26371 ( n16040 , n13353 , n3257 );
    not g26372 ( n19614 , n14160 );
    or g26373 ( n29940 , n15488 , n20290 );
    not g26374 ( n31994 , n23187 );
    xnor g26375 ( n17646 , n15999 , n7414 );
    or g26376 ( n14651 , n27728 , n31684 );
    and g26377 ( n7693 , n609 , n5842 );
    and g26378 ( n24497 , n2455 , n25327 );
    or g26379 ( n4028 , n21899 , n16320 );
    and g26380 ( n20777 , n21792 , n10491 );
    and g26381 ( n17845 , n9134 , n8370 );
    not g26382 ( n13903 , n11518 );
    nor g26383 ( n29215 , n16633 , n2116 );
    and g26384 ( n926 , n6822 , n19221 );
    and g26385 ( n6733 , n4936 , n1291 );
    xnor g26386 ( n19752 , n8442 , n6660 );
    or g26387 ( n14435 , n2138 , n16555 );
    nor g26388 ( n6329 , n29447 , n25689 );
    and g26389 ( n15462 , n8600 , n17331 );
    or g26390 ( n26015 , n6212 , n25060 );
    or g26391 ( n4770 , n25219 , n2416 );
    or g26392 ( n28708 , n31183 , n29419 );
    not g26393 ( n29826 , n20569 );
    not g26394 ( n385 , n9543 );
    or g26395 ( n25865 , n9509 , n4517 );
    xnor g26396 ( n30898 , n8887 , n21334 );
    or g26397 ( n26223 , n4118 , n24263 );
    not g26398 ( n6117 , n29930 );
    xnor g26399 ( n13048 , n1816 , n16485 );
    not g26400 ( n27482 , n7129 );
    xor g26401 ( n18184 , n25464 , n11866 );
    and g26402 ( n29313 , n7498 , n25258 );
    xnor g26403 ( n1638 , n13664 , n21067 );
    not g26404 ( n5995 , n17132 );
    or g26405 ( n30661 , n18071 , n21417 );
    and g26406 ( n27666 , n29428 , n18813 );
    and g26407 ( n21330 , n27835 , n6265 );
    or g26408 ( n2284 , n9281 , n21091 );
    xnor g26409 ( n22863 , n90 , n15413 );
    nor g26410 ( n22446 , n28110 , n23184 );
    nor g26411 ( n14342 , n31839 , n25372 );
    xnor g26412 ( n9443 , n12112 , n22837 );
    and g26413 ( n14801 , n31275 , n21699 );
    or g26414 ( n21983 , n25534 , n23990 );
    or g26415 ( n17907 , n6901 , n4936 );
    not g26416 ( n11747 , n30126 );
    and g26417 ( n15202 , n578 , n1927 );
    or g26418 ( n25722 , n26636 , n11998 );
    or g26419 ( n16750 , n11195 , n7546 );
    or g26420 ( n3974 , n13186 , n1807 );
    xnor g26421 ( n19610 , n28357 , n244 );
    and g26422 ( n19688 , n11011 , n5138 );
    and g26423 ( n30833 , n20081 , n13108 );
    not g26424 ( n24897 , n9596 );
    and g26425 ( n27336 , n25326 , n31635 );
    xnor g26426 ( n14397 , n13828 , n28040 );
    not g26427 ( n2107 , n12640 );
    or g26428 ( n21747 , n2765 , n9022 );
    and g26429 ( n4896 , n23451 , n31823 );
    xor g26430 ( n25121 , n26916 , n26824 );
    not g26431 ( n27357 , n5205 );
    xnor g26432 ( n31818 , n21341 , n12306 );
    not g26433 ( n23777 , n23419 );
    xnor g26434 ( n27456 , n24992 , n25053 );
    xor g26435 ( n19574 , n8368 , n21231 );
    and g26436 ( n20172 , n7275 , n29694 );
    not g26437 ( n11008 , n20349 );
    nor g26438 ( n10942 , n13478 , n12214 );
    nor g26439 ( n24298 , n31502 , n3491 );
    or g26440 ( n17409 , n21064 , n11950 );
    and g26441 ( n17836 , n4454 , n24787 );
    and g26442 ( n4016 , n29654 , n16688 );
    nor g26443 ( n30953 , n19701 , n10911 );
    nor g26444 ( n29428 , n30422 , n28186 );
    and g26445 ( n26303 , n15455 , n484 );
    not g26446 ( n13040 , n4996 );
    xnor g26447 ( n13551 , n23820 , n7768 );
    or g26448 ( n18481 , n834 , n16616 );
    and g26449 ( n11857 , n815 , n6785 );
    and g26450 ( n2579 , n30877 , n3652 );
    xor g26451 ( n15039 , n12603 , n1693 );
    or g26452 ( n18021 , n23754 , n4029 );
    nor g26453 ( n28304 , n24178 , n2051 );
    nor g26454 ( n21473 , n5113 , n10569 );
    xnor g26455 ( n17396 , n15741 , n11995 );
    and g26456 ( n3562 , n28928 , n30439 );
    xnor g26457 ( n29910 , n22662 , n9605 );
    and g26458 ( n26652 , n21012 , n1152 );
    or g26459 ( n28977 , n15549 , n5040 );
    or g26460 ( n9156 , n3487 , n20204 );
    or g26461 ( n19065 , n2050 , n6845 );
    not g26462 ( n11109 , n29233 );
    nor g26463 ( n2134 , n8337 , n29865 );
    not g26464 ( n13697 , n19358 );
    or g26465 ( n1110 , n10036 , n2295 );
    not g26466 ( n17027 , n7453 );
    xnor g26467 ( n17250 , n10810 , n11305 );
    not g26468 ( n17878 , n6783 );
    nor g26469 ( n10112 , n20198 , n20490 );
    xnor g26470 ( n13121 , n11587 , n15266 );
    or g26471 ( n23612 , n10732 , n12463 );
    xnor g26472 ( n7019 , n12312 , n10737 );
    not g26473 ( n27695 , n20495 );
    and g26474 ( n31451 , n5398 , n3132 );
    nor g26475 ( n17212 , n28177 , n25541 );
    xnor g26476 ( n15155 , n17565 , n476 );
    xnor g26477 ( n31740 , n7234 , n9469 );
    not g26478 ( n20574 , n29407 );
    nor g26479 ( n25861 , n19300 , n18746 );
    and g26480 ( n27382 , n491 , n25888 );
    xnor g26481 ( n26674 , n22819 , n4375 );
    not g26482 ( n5415 , n16001 );
    xnor g26483 ( n14383 , n6492 , n14037 );
    not g26484 ( n24104 , n16881 );
    xnor g26485 ( n25095 , n30639 , n21261 );
    and g26486 ( n16474 , n30276 , n8133 );
    or g26487 ( n29048 , n20155 , n31817 );
    nor g26488 ( n14460 , n12104 , n12614 );
    not g26489 ( n23003 , n6448 );
    xnor g26490 ( n14825 , n24159 , n19970 );
    not g26491 ( n28165 , n29435 );
    xnor g26492 ( n9439 , n30370 , n3163 );
    nor g26493 ( n24963 , n6372 , n29320 );
    and g26494 ( n29743 , n30715 , n16631 );
    or g26495 ( n1619 , n23590 , n24031 );
    xnor g26496 ( n29023 , n6752 , n565 );
    xnor g26497 ( n18015 , n13797 , n30245 );
    nor g26498 ( n857 , n13656 , n512 );
    or g26499 ( n27665 , n495 , n3343 );
    not g26500 ( n21241 , n2485 );
    not g26501 ( n15526 , n23341 );
    not g26502 ( n244 , n4928 );
    not g26503 ( n13220 , n10959 );
    xnor g26504 ( n1961 , n16154 , n13737 );
    and g26505 ( n23161 , n16632 , n16543 );
    not g26506 ( n25237 , n4796 );
    xnor g26507 ( n13906 , n26082 , n25793 );
    and g26508 ( n22987 , n10273 , n9305 );
    xnor g26509 ( n2006 , n14585 , n23943 );
    or g26510 ( n14879 , n3005 , n30144 );
    xnor g26511 ( n24181 , n19994 , n18374 );
    xnor g26512 ( n16054 , n3586 , n10965 );
    nor g26513 ( n14019 , n19220 , n19622 );
    not g26514 ( n30602 , n4601 );
    and g26515 ( n23719 , n17507 , n28140 );
    xnor g26516 ( n20346 , n11257 , n17617 );
    xor g26517 ( n28667 , n12471 , n9604 );
    xor g26518 ( n28278 , n9925 , n74 );
    or g26519 ( n25640 , n28700 , n13523 );
    not g26520 ( n17704 , n1439 );
    xnor g26521 ( n26011 , n5522 , n27407 );
    and g26522 ( n9557 , n30857 , n24380 );
    or g26523 ( n26041 , n2176 , n21995 );
    xnor g26524 ( n5866 , n23849 , n1405 );
    xnor g26525 ( n17713 , n23066 , n943 );
    xnor g26526 ( n5133 , n17189 , n6699 );
    xnor g26527 ( n26741 , n8312 , n27630 );
    not g26528 ( n20611 , n6076 );
    not g26529 ( n16028 , n24929 );
    or g26530 ( n12424 , n30130 , n2089 );
    not g26531 ( n28408 , n21216 );
    nor g26532 ( n16805 , n8321 , n7209 );
    xnor g26533 ( n31066 , n31532 , n30968 );
    or g26534 ( n11650 , n23817 , n6818 );
    nor g26535 ( n17445 , n22421 , n29109 );
    not g26536 ( n4188 , n19494 );
    not g26537 ( n2160 , n13067 );
    or g26538 ( n18574 , n3836 , n20696 );
    not g26539 ( n12159 , n30186 );
    xnor g26540 ( n21246 , n23031 , n14065 );
    and g26541 ( n27137 , n8537 , n2752 );
    not g26542 ( n19582 , n28267 );
    not g26543 ( n15547 , n9138 );
    buf g26544 ( n9638 , n25460 );
    and g26545 ( n20969 , n6008 , n10819 );
    and g26546 ( n6242 , n28659 , n30157 );
    not g26547 ( n24608 , n15971 );
    xnor g26548 ( n9613 , n5597 , n25614 );
    and g26549 ( n25029 , n16596 , n10258 );
    xnor g26550 ( n21340 , n30866 , n8321 );
    or g26551 ( n24501 , n25477 , n1661 );
    or g26552 ( n13297 , n23462 , n1158 );
    xnor g26553 ( n15820 , n21993 , n23306 );
    xnor g26554 ( n24389 , n5060 , n9163 );
    not g26555 ( n7010 , n14960 );
    or g26556 ( n24045 , n20195 , n7841 );
    and g26557 ( n28516 , n27545 , n6450 );
    not g26558 ( n14848 , n24736 );
    and g26559 ( n20414 , n31239 , n19138 );
    and g26560 ( n28540 , n31712 , n28534 );
    or g26561 ( n31039 , n29133 , n15646 );
    xnor g26562 ( n14788 , n19068 , n3426 );
    and g26563 ( n1563 , n21441 , n21963 );
    xor g26564 ( n15162 , n23722 , n21620 );
    or g26565 ( n2140 , n14172 , n13107 );
    nor g26566 ( n12290 , n3275 , n8334 );
    xnor g26567 ( n14034 , n22457 , n22089 );
    not g26568 ( n6425 , n22816 );
    xnor g26569 ( n20002 , n23683 , n3916 );
    and g26570 ( n1443 , n28792 , n21608 );
    or g26571 ( n8690 , n1980 , n11950 );
    or g26572 ( n6079 , n17617 , n1817 );
    xnor g26573 ( n16706 , n23878 , n7198 );
    xnor g26574 ( n7605 , n5387 , n6295 );
    xnor g26575 ( n9311 , n31262 , n3274 );
    or g26576 ( n20001 , n26856 , n2976 );
    xnor g26577 ( n17038 , n512 , n30455 );
    or g26578 ( n879 , n12083 , n8858 );
    and g26579 ( n26118 , n21038 , n18394 );
    or g26580 ( n4400 , n17138 , n12778 );
    and g26581 ( n12637 , n29371 , n26224 );
    and g26582 ( n26927 , n31025 , n26253 );
    not g26583 ( n4332 , n375 );
    xnor g26584 ( n22600 , n281 , n6616 );
    nor g26585 ( n20222 , n29243 , n22531 );
    or g26586 ( n10919 , n7651 , n20107 );
    xnor g26587 ( n24753 , n25481 , n23057 );
    xnor g26588 ( n4504 , n7670 , n27443 );
    nor g26589 ( n23986 , n30882 , n265 );
    or g26590 ( n13997 , n27911 , n22147 );
    nor g26591 ( n3487 , n26489 , n25280 );
    nor g26592 ( n24679 , n14503 , n31420 );
    xnor g26593 ( n23749 , n3851 , n396 );
    and g26594 ( n28672 , n9931 , n19960 );
    not g26595 ( n1203 , n25206 );
    not g26596 ( n29854 , n28571 );
    not g26597 ( n11646 , n20515 );
    not g26598 ( n10302 , n9835 );
    xnor g26599 ( n22681 , n19062 , n20198 );
    or g26600 ( n28726 , n15873 , n5596 );
    not g26601 ( n28331 , n17263 );
    not g26602 ( n31676 , n10334 );
    nor g26603 ( n20751 , n1141 , n11447 );
    not g26604 ( n4898 , n27184 );
    or g26605 ( n14379 , n22665 , n15036 );
    and g26606 ( n27582 , n17778 , n6888 );
    or g26607 ( n21965 , n17008 , n15045 );
    xnor g26608 ( n2911 , n22004 , n24441 );
    or g26609 ( n30060 , n30525 , n29632 );
    buf g26610 ( n9396 , n19137 );
    xnor g26611 ( n31619 , n20953 , n21454 );
    xnor g26612 ( n17712 , n1211 , n25665 );
    xnor g26613 ( n19771 , n15009 , n16019 );
    xnor g26614 ( n17773 , n9910 , n26345 );
    not g26615 ( n29255 , n110 );
    or g26616 ( n20511 , n14291 , n23192 );
    or g26617 ( n24232 , n16283 , n18580 );
    or g26618 ( n25919 , n5880 , n25620 );
    and g26619 ( n24982 , n24470 , n30743 );
    or g26620 ( n15269 , n23040 , n11439 );
    and g26621 ( n28371 , n27038 , n19576 );
    not g26622 ( n8816 , n1995 );
    not g26623 ( n31222 , n31653 );
    xor g26624 ( n27963 , n26350 , n16822 );
    xnor g26625 ( n17687 , n17584 , n10713 );
    not g26626 ( n25721 , n8191 );
    and g26627 ( n29834 , n23296 , n14596 );
    and g26628 ( n21198 , n7402 , n22096 );
    nor g26629 ( n21847 , n11870 , n11363 );
    not g26630 ( n12087 , n12641 );
    xnor g26631 ( n12862 , n2294 , n31426 );
    and g26632 ( n7298 , n8203 , n9988 );
    not g26633 ( n19420 , n3022 );
    not g26634 ( n22868 , n8289 );
    xor g26635 ( n23769 , n13443 , n17526 );
    and g26636 ( n4477 , n1379 , n16105 );
    xnor g26637 ( n20953 , n23812 , n25382 );
    and g26638 ( n24898 , n4101 , n25850 );
    or g26639 ( n506 , n15563 , n29998 );
    or g26640 ( n26618 , n29586 , n15540 );
    or g26641 ( n28897 , n15281 , n29618 );
    or g26642 ( n12381 , n16673 , n15218 );
    xnor g26643 ( n5475 , n386 , n7315 );
    xnor g26644 ( n17291 , n19605 , n21865 );
    or g26645 ( n27540 , n30167 , n7391 );
    and g26646 ( n25928 , n19850 , n25785 );
    xnor g26647 ( n8385 , n26440 , n26684 );
    not g26648 ( n17262 , n5496 );
    or g26649 ( n20422 , n1331 , n1865 );
    and g26650 ( n11571 , n123 , n18495 );
    and g26651 ( n21240 , n1905 , n16510 );
    and g26652 ( n20153 , n5845 , n26210 );
    or g26653 ( n28876 , n13035 , n13193 );
    xnor g26654 ( n20749 , n31441 , n4405 );
    or g26655 ( n17962 , n326 , n15925 );
    not g26656 ( n29896 , n12725 );
    and g26657 ( n1140 , n20984 , n5508 );
    xnor g26658 ( n26348 , n31414 , n18253 );
    xnor g26659 ( n19537 , n29852 , n19904 );
    nor g26660 ( n7944 , n5041 , n20397 );
    not g26661 ( n10947 , n11222 );
    not g26662 ( n24437 , n25000 );
    xnor g26663 ( n21639 , n30262 , n31326 );
    xnor g26664 ( n9130 , n713 , n26191 );
    not g26665 ( n14201 , n17990 );
    xnor g26666 ( n4032 , n2692 , n1365 );
    and g26667 ( n13926 , n14953 , n15630 );
    or g26668 ( n28339 , n28990 , n1797 );
    not g26669 ( n13712 , n9113 );
    not g26670 ( n18558 , n18203 );
    not g26671 ( n8505 , n6824 );
    and g26672 ( n25114 , n27823 , n12272 );
    xnor g26673 ( n14745 , n22678 , n13410 );
    not g26674 ( n29336 , n3700 );
    xnor g26675 ( n14044 , n13471 , n5317 );
    xnor g26676 ( n23869 , n22318 , n6250 );
    xnor g26677 ( n13299 , n23444 , n2146 );
    nor g26678 ( n22030 , n11218 , n2447 );
    xnor g26679 ( n23187 , n27463 , n6729 );
    or g26680 ( n6688 , n26735 , n2990 );
    and g26681 ( n758 , n15228 , n30458 );
    not g26682 ( n28376 , n30805 );
    not g26683 ( n16794 , n863 );
    or g26684 ( n22108 , n22911 , n373 );
    or g26685 ( n30960 , n14792 , n20633 );
    xnor g26686 ( n19379 , n9011 , n21186 );
    and g26687 ( n31151 , n717 , n22069 );
    nor g26688 ( n5161 , n20748 , n9540 );
    nor g26689 ( n20184 , n12298 , n27271 );
    nor g26690 ( n29331 , n16799 , n18135 );
    and g26691 ( n26406 , n10952 , n30594 );
    or g26692 ( n29352 , n4811 , n17631 );
    and g26693 ( n5726 , n30437 , n28888 );
    xnor g26694 ( n11938 , n21927 , n19188 );
    or g26695 ( n5843 , n25546 , n4176 );
    not g26696 ( n17611 , n12625 );
    nor g26697 ( n28149 , n7767 , n25982 );
    not g26698 ( n8269 , n18184 );
    and g26699 ( n13578 , n27346 , n19533 );
    or g26700 ( n20068 , n13160 , n22127 );
    and g26701 ( n20757 , n4866 , n4782 );
    or g26702 ( n18978 , n6324 , n24923 );
    xnor g26703 ( n6579 , n4721 , n18758 );
    and g26704 ( n10779 , n24876 , n21322 );
    or g26705 ( n5844 , n25884 , n7469 );
    nor g26706 ( n10453 , n18735 , n27411 );
    or g26707 ( n14188 , n2444 , n4185 );
    not g26708 ( n7996 , n11964 );
    or g26709 ( n3729 , n3508 , n17977 );
    xnor g26710 ( n1084 , n18428 , n904 );
    xnor g26711 ( n2626 , n1171 , n8927 );
    or g26712 ( n2013 , n21150 , n723 );
    not g26713 ( n1606 , n6599 );
    and g26714 ( n27036 , n7189 , n6513 );
    not g26715 ( n20639 , n3849 );
    not g26716 ( n15391 , n23833 );
    not g26717 ( n30699 , n21476 );
    xnor g26718 ( n24617 , n1428 , n25660 );
    not g26719 ( n10534 , n8620 );
    or g26720 ( n10161 , n28953 , n22082 );
    not g26721 ( n516 , n14112 );
    or g26722 ( n4385 , n22900 , n4699 );
    not g26723 ( n8367 , n7159 );
    xnor g26724 ( n26517 , n546 , n27503 );
    xnor g26725 ( n1228 , n11526 , n2603 );
    or g26726 ( n1071 , n11253 , n12193 );
    not g26727 ( n15648 , n31019 );
    or g26728 ( n25155 , n20395 , n1914 );
    not g26729 ( n5825 , n11206 );
    not g26730 ( n15424 , n1039 );
    and g26731 ( n18532 , n30104 , n8549 );
    or g26732 ( n22293 , n25017 , n4766 );
    xnor g26733 ( n31544 , n16031 , n24436 );
    xnor g26734 ( n3290 , n4370 , n26208 );
    not g26735 ( n12226 , n26378 );
    xnor g26736 ( n8605 , n7731 , n15512 );
    or g26737 ( n21894 , n17995 , n4815 );
    nor g26738 ( n384 , n30792 , n30352 );
    xnor g26739 ( n22652 , n13339 , n17955 );
    nor g26740 ( n22895 , n1499 , n528 );
    xnor g26741 ( n10403 , n11400 , n12216 );
    nor g26742 ( n31284 , n14411 , n29847 );
    buf g26743 ( n8577 , n11756 );
    and g26744 ( n1782 , n24045 , n27240 );
    not g26745 ( n1566 , n27366 );
    nor g26746 ( n1626 , n30290 , n7280 );
    or g26747 ( n14278 , n837 , n6090 );
    or g26748 ( n19520 , n25070 , n2793 );
    xnor g26749 ( n15658 , n17045 , n8508 );
    not g26750 ( n2082 , n1934 );
    not g26751 ( n23669 , n23577 );
    or g26752 ( n954 , n5233 , n19966 );
    xnor g26753 ( n12090 , n26458 , n24563 );
    nor g26754 ( n22912 , n21136 , n18551 );
    not g26755 ( n3693 , n1971 );
    xnor g26756 ( n23189 , n14115 , n23507 );
    xnor g26757 ( n26440 , n11081 , n22243 );
    and g26758 ( n27264 , n29903 , n5282 );
    or g26759 ( n6513 , n15382 , n4174 );
    xnor g26760 ( n20224 , n22420 , n30022 );
    nor g26761 ( n2518 , n256 , n331 );
    nor g26762 ( n10311 , n14477 , n27411 );
    not g26763 ( n7781 , n15298 );
    not g26764 ( n13120 , n19428 );
    not g26765 ( n5483 , n3996 );
    nor g26766 ( n19257 , n25179 , n17126 );
    not g26767 ( n28403 , n24569 );
    xnor g26768 ( n13962 , n18788 , n26029 );
    not g26769 ( n9538 , n25760 );
    or g26770 ( n24654 , n9286 , n8987 );
    not g26771 ( n29371 , n10859 );
    not g26772 ( n1702 , n11938 );
    not g26773 ( n10347 , n11616 );
    or g26774 ( n28014 , n18999 , n1341 );
    and g26775 ( n3463 , n3797 , n20487 );
    not g26776 ( n7284 , n24769 );
    not g26777 ( n13062 , n22622 );
    xnor g26778 ( n19625 , n9542 , n27935 );
    xnor g26779 ( n15833 , n15889 , n28305 );
    xnor g26780 ( n18284 , n25114 , n3657 );
    not g26781 ( n5118 , n1557 );
    xnor g26782 ( n11565 , n14091 , n25798 );
    xnor g26783 ( n23764 , n1780 , n20394 );
    or g26784 ( n24632 , n24320 , n23606 );
    and g26785 ( n22725 , n18991 , n30267 );
    xnor g26786 ( n9487 , n18551 , n15749 );
    not g26787 ( n19710 , n30863 );
    or g26788 ( n17451 , n5948 , n23202 );
    or g26789 ( n27702 , n31920 , n30751 );
    nor g26790 ( n604 , n16799 , n21720 );
    or g26791 ( n20094 , n7465 , n3991 );
    xnor g26792 ( n3394 , n7952 , n3746 );
    xnor g26793 ( n27178 , n17854 , n6633 );
    or g26794 ( n5124 , n16526 , n15412 );
    xnor g26795 ( n21315 , n30887 , n23960 );
    not g26796 ( n3073 , n16266 );
    xnor g26797 ( n19662 , n13527 , n24524 );
    or g26798 ( n15028 , n23349 , n23258 );
    or g26799 ( n14165 , n3136 , n21144 );
    or g26800 ( n13231 , n27307 , n16923 );
    not g26801 ( n17000 , n13044 );
    not g26802 ( n26204 , n14598 );
    not g26803 ( n28999 , n22531 );
    or g26804 ( n25258 , n14792 , n22569 );
    or g26805 ( n17590 , n20135 , n12372 );
    xnor g26806 ( n14262 , n21695 , n13438 );
    not g26807 ( n5064 , n29474 );
    and g26808 ( n27312 , n27563 , n31565 );
    not g26809 ( n14982 , n5345 );
    xnor g26810 ( n26375 , n28829 , n20390 );
    nor g26811 ( n15205 , n18247 , n890 );
    not g26812 ( n27954 , n28448 );
    not g26813 ( n21819 , n25495 );
    xnor g26814 ( n14273 , n12073 , n24132 );
    nor g26815 ( n1400 , n6086 , n6168 );
    or g26816 ( n21794 , n2411 , n10007 );
    xnor g26817 ( n31883 , n24784 , n17019 );
    and g26818 ( n26629 , n30258 , n8008 );
    xnor g26819 ( n9474 , n6474 , n26191 );
    or g26820 ( n5140 , n14557 , n13939 );
    or g26821 ( n633 , n20647 , n26119 );
    or g26822 ( n586 , n31770 , n1674 );
    or g26823 ( n26876 , n31281 , n27055 );
    not g26824 ( n8268 , n24113 );
    or g26825 ( n19914 , n28701 , n8437 );
    and g26826 ( n23604 , n23665 , n11546 );
    xnor g26827 ( n22814 , n3969 , n17234 );
    xnor g26828 ( n16210 , n1720 , n29249 );
    or g26829 ( n28443 , n31345 , n11952 );
    not g26830 ( n22208 , n4052 );
    and g26831 ( n20220 , n18668 , n22045 );
    or g26832 ( n9307 , n17417 , n16898 );
    xnor g26833 ( n2303 , n24328 , n7278 );
    not g26834 ( n21863 , n9743 );
    buf g26835 ( n25856 , n11896 );
    not g26836 ( n11912 , n11552 );
    not g26837 ( n13476 , n20210 );
    and g26838 ( n15134 , n21794 , n13127 );
    or g26839 ( n13165 , n19401 , n7020 );
    or g26840 ( n30478 , n2778 , n24637 );
    nor g26841 ( n24033 , n4987 , n28144 );
    not g26842 ( n29950 , n9525 );
    and g26843 ( n28644 , n3367 , n11984 );
    xnor g26844 ( n949 , n8846 , n26055 );
    or g26845 ( n20065 , n478 , n21336 );
    xnor g26846 ( n15438 , n13558 , n5230 );
    xnor g26847 ( n31124 , n20408 , n12668 );
    not g26848 ( n10812 , n29905 );
    nor g26849 ( n5771 , n11345 , n2020 );
    xnor g26850 ( n26197 , n26142 , n11185 );
    not g26851 ( n10881 , n8251 );
    or g26852 ( n28764 , n20995 , n15641 );
    xnor g26853 ( n31058 , n27862 , n23806 );
    xnor g26854 ( n9545 , n3898 , n29510 );
    xnor g26855 ( n31261 , n11426 , n21963 );
    not g26856 ( n9824 , n10145 );
    not g26857 ( n7424 , n3701 );
    nor g26858 ( n30052 , n6637 , n26549 );
    xnor g26859 ( n19925 , n5325 , n1059 );
    not g26860 ( n7558 , n7330 );
    and g26861 ( n1069 , n10768 , n14573 );
    not g26862 ( n780 , n22395 );
    and g26863 ( n7515 , n15042 , n13784 );
    xnor g26864 ( n20952 , n16214 , n8145 );
    and g26865 ( n31685 , n25376 , n30310 );
    xnor g26866 ( n25112 , n2260 , n16365 );
    or g26867 ( n21861 , n10991 , n12093 );
    or g26868 ( n11111 , n26096 , n8212 );
    xnor g26869 ( n22617 , n9506 , n725 );
    and g26870 ( n7253 , n19268 , n6926 );
    nor g26871 ( n22035 , n5327 , n2877 );
    xor g26872 ( n25415 , n16188 , n23373 );
    or g26873 ( n25705 , n30485 , n16296 );
    not g26874 ( n1319 , n14867 );
    not g26875 ( n23056 , n2443 );
    and g26876 ( n161 , n13513 , n24329 );
    not g26877 ( n4909 , n15696 );
    xnor g26878 ( n31625 , n28190 , n21303 );
    or g26879 ( n27547 , n10458 , n21513 );
    or g26880 ( n1657 , n14553 , n6473 );
    xnor g26881 ( n20237 , n9852 , n11197 );
    not g26882 ( n18884 , n8232 );
    not g26883 ( n9300 , n14779 );
    xnor g26884 ( n27801 , n23271 , n29108 );
    not g26885 ( n31759 , n8266 );
    and g26886 ( n26076 , n6702 , n27699 );
    or g26887 ( n3685 , n5408 , n19012 );
    and g26888 ( n581 , n23782 , n6922 );
    xnor g26889 ( n29583 , n16286 , n3713 );
    or g26890 ( n2276 , n5032 , n15128 );
    not g26891 ( n12970 , n12607 );
    or g26892 ( n22465 , n312 , n678 );
    xnor g26893 ( n9524 , n14090 , n15588 );
    xnor g26894 ( n18400 , n19000 , n12971 );
    xnor g26895 ( n3480 , n11582 , n17312 );
    not g26896 ( n15689 , n30894 );
    nor g26897 ( n17239 , n24988 , n3210 );
    or g26898 ( n11006 , n17441 , n11063 );
    and g26899 ( n3757 , n12162 , n2604 );
    and g26900 ( n25377 , n3623 , n15905 );
    not g26901 ( n15078 , n3239 );
    or g26902 ( n27035 , n8001 , n19325 );
    not g26903 ( n24069 , n6740 );
    xnor g26904 ( n8479 , n31697 , n27071 );
    xnor g26905 ( n18686 , n8221 , n6694 );
    and g26906 ( n1243 , n23200 , n5259 );
    xnor g26907 ( n31603 , n26288 , n11388 );
    xnor g26908 ( n16783 , n15765 , n23280 );
    nor g26909 ( n5603 , n20799 , n2939 );
    not g26910 ( n18530 , n28729 );
    xnor g26911 ( n7264 , n5984 , n11132 );
    or g26912 ( n21155 , n13418 , n10009 );
    xnor g26913 ( n24283 , n11821 , n26698 );
    or g26914 ( n9459 , n27948 , n19678 );
    xor g26915 ( n1557 , n9457 , n2726 );
    not g26916 ( n13312 , n810 );
    xnor g26917 ( n5109 , n21499 , n27753 );
    xnor g26918 ( n20180 , n30043 , n11908 );
    or g26919 ( n10513 , n29952 , n20775 );
    xnor g26920 ( n6811 , n20674 , n19880 );
    or g26921 ( n11224 , n16518 , n26184 );
    nor g26922 ( n11019 , n7593 , n29751 );
    not g26923 ( n16793 , n4952 );
    xnor g26924 ( n16249 , n30125 , n11627 );
    nor g26925 ( n4961 , n11920 , n11943 );
    not g26926 ( n24212 , n5328 );
    xnor g26927 ( n17780 , n5934 , n22946 );
    or g26928 ( n14436 , n979 , n9346 );
    and g26929 ( n30763 , n11432 , n11480 );
    xnor g26930 ( n12117 , n24270 , n6902 );
    and g26931 ( n27118 , n18562 , n22550 );
    xnor g26932 ( n12509 , n9080 , n16273 );
    and g26933 ( n17431 , n18597 , n9606 );
    or g26934 ( n19455 , n19943 , n15452 );
    or g26935 ( n31527 , n445 , n18389 );
    not g26936 ( n11798 , n19496 );
    and g26937 ( n28119 , n14138 , n17668 );
    and g26938 ( n12456 , n9856 , n13987 );
    nor g26939 ( n26366 , n10202 , n4032 );
    xnor g26940 ( n21422 , n5790 , n15839 );
    not g26941 ( n1649 , n12279 );
    nor g26942 ( n30272 , n19720 , n15557 );
    xor g26943 ( n7928 , n23899 , n27057 );
    and g26944 ( n5504 , n26506 , n28753 );
    not g26945 ( n27866 , n5089 );
    or g26946 ( n20910 , n3485 , n4393 );
    xnor g26947 ( n8074 , n5798 , n18613 );
    and g26948 ( n2973 , n9960 , n17648 );
    not g26949 ( n7587 , n30479 );
    nor g26950 ( n26342 , n17755 , n5833 );
    or g26951 ( n9238 , n2736 , n26458 );
    xnor g26952 ( n22447 , n19367 , n15380 );
    and g26953 ( n7769 , n29537 , n26154 );
    or g26954 ( n20892 , n20773 , n1631 );
    not g26955 ( n20040 , n22516 );
    xnor g26956 ( n15759 , n9247 , n31647 );
    or g26957 ( n26714 , n433 , n30878 );
    xnor g26958 ( n27365 , n14681 , n7111 );
    and g26959 ( n1693 , n18136 , n3342 );
    xnor g26960 ( n16597 , n29163 , n10713 );
    not g26961 ( n8446 , n28638 );
    not g26962 ( n18327 , n26989 );
    xor g26963 ( n8004 , n2794 , n26887 );
    or g26964 ( n8843 , n16895 , n21601 );
    not g26965 ( n9962 , n9653 );
    not g26966 ( n29411 , n28562 );
    nor g26967 ( n15606 , n25856 , n12971 );
    nor g26968 ( n1493 , n29008 , n26991 );
    or g26969 ( n4401 , n9123 , n14614 );
    not g26970 ( n2956 , n28766 );
    or g26971 ( n17507 , n29442 , n24044 );
    and g26972 ( n25681 , n6835 , n22658 );
    not g26973 ( n4483 , n17173 );
    nor g26974 ( n24838 , n3668 , n20021 );
    not g26975 ( n23495 , n27359 );
    xnor g26976 ( n28956 , n30190 , n1042 );
    xnor g26977 ( n2205 , n17369 , n22013 );
    or g26978 ( n30011 , n22512 , n16779 );
    or g26979 ( n4794 , n23209 , n31288 );
    xnor g26980 ( n4697 , n7378 , n20365 );
    and g26981 ( n30023 , n14694 , n16815 );
    not g26982 ( n7872 , n22413 );
    not g26983 ( n22759 , n588 );
    not g26984 ( n15698 , n21068 );
    xnor g26985 ( n25936 , n24451 , n29702 );
    xnor g26986 ( n20121 , n10683 , n7800 );
    not g26987 ( n25344 , n20819 );
    xnor g26988 ( n25020 , n5866 , n3563 );
    xnor g26989 ( n11068 , n14974 , n757 );
    or g26990 ( n26136 , n6439 , n4320 );
    not g26991 ( n9807 , n6456 );
    nor g26992 ( n16379 , n31975 , n29557 );
    not g26993 ( n22318 , n15190 );
    and g26994 ( n6255 , n21108 , n29205 );
    or g26995 ( n28251 , n20561 , n26587 );
    not g26996 ( n3545 , n13712 );
    not g26997 ( n10169 , n10404 );
    xnor g26998 ( n20022 , n25252 , n14925 );
    not g26999 ( n17615 , n8782 );
    not g27000 ( n28601 , n4384 );
    and g27001 ( n22781 , n26201 , n7802 );
    not g27002 ( n27360 , n19525 );
    and g27003 ( n1846 , n3862 , n11007 );
    not g27004 ( n3388 , n31391 );
    not g27005 ( n31866 , n19896 );
    or g27006 ( n11214 , n17326 , n21416 );
    and g27007 ( n14108 , n11290 , n24350 );
    not g27008 ( n16465 , n18840 );
    or g27009 ( n21486 , n2963 , n27250 );
    xnor g27010 ( n24087 , n14643 , n17674 );
    xnor g27011 ( n20602 , n17097 , n122 );
    and g27012 ( n10046 , n781 , n10581 );
    or g27013 ( n8366 , n19742 , n4010 );
    not g27014 ( n25351 , n7980 );
    xor g27015 ( n11618 , n1589 , n30297 );
    or g27016 ( n17625 , n23254 , n8760 );
    not g27017 ( n1680 , n20954 );
    or g27018 ( n31746 , n12055 , n7496 );
    not g27019 ( n13649 , n25637 );
    and g27020 ( n21784 , n16514 , n29552 );
    not g27021 ( n14307 , n17953 );
    or g27022 ( n2365 , n11980 , n19751 );
    or g27023 ( n7660 , n28402 , n21482 );
    not g27024 ( n150 , n23306 );
    not g27025 ( n2693 , n7925 );
    or g27026 ( n10191 , n4224 , n10281 );
    or g27027 ( n6802 , n24978 , n30237 );
    and g27028 ( n917 , n11790 , n4005 );
    not g27029 ( n9213 , n27967 );
    not g27030 ( n10066 , n977 );
    xnor g27031 ( n5405 , n10770 , n23281 );
    not g27032 ( n29239 , n988 );
    nor g27033 ( n19944 , n109 , n18807 );
    or g27034 ( n19807 , n20558 , n16879 );
    nor g27035 ( n14086 , n10044 , n4663 );
    not g27036 ( n8117 , n25198 );
    not g27037 ( n12187 , n4568 );
    or g27038 ( n12761 , n25532 , n18496 );
    xnor g27039 ( n10781 , n3056 , n32009 );
    xnor g27040 ( n24588 , n26114 , n4836 );
    not g27041 ( n5432 , n10467 );
    xnor g27042 ( n25460 , n22639 , n1974 );
    not g27043 ( n30108 , n17477 );
    xnor g27044 ( n10975 , n851 , n19384 );
    xor g27045 ( n3808 , n9307 , n10949 );
    xnor g27046 ( n24714 , n23097 , n15999 );
    or g27047 ( n7946 , n12961 , n22547 );
    or g27048 ( n6023 , n24787 , n1956 );
    xnor g27049 ( n9064 , n17089 , n22422 );
    not g27050 ( n17831 , n26689 );
    not g27051 ( n29808 , n15940 );
    not g27052 ( n8345 , n26695 );
    or g27053 ( n9295 , n22596 , n18420 );
    or g27054 ( n941 , n27605 , n14000 );
    nor g27055 ( n6326 , n28368 , n15669 );
    xnor g27056 ( n29119 , n19020 , n13520 );
    or g27057 ( n224 , n23577 , n18529 );
    xnor g27058 ( n19934 , n13297 , n27750 );
    or g27059 ( n31167 , n14878 , n27796 );
    not g27060 ( n3173 , n14816 );
    xnor g27061 ( n24451 , n12143 , n22866 );
    and g27062 ( n3672 , n4281 , n10505 );
    xnor g27063 ( n31343 , n6605 , n1525 );
    not g27064 ( n20118 , n9043 );
    xor g27065 ( n25476 , n24980 , n20435 );
    xnor g27066 ( n8347 , n7814 , n15634 );
    not g27067 ( n17350 , n7462 );
    nor g27068 ( n23110 , n14604 , n6613 );
    not g27069 ( n11838 , n30233 );
    xnor g27070 ( n26957 , n26952 , n26461 );
    xor g27071 ( n29389 , n21859 , n15570 );
    and g27072 ( n2119 , n18194 , n18376 );
    or g27073 ( n10650 , n13040 , n28346 );
    or g27074 ( n15229 , n25089 , n30552 );
    and g27075 ( n6654 , n30140 , n9622 );
    nor g27076 ( n17940 , n4686 , n15838 );
    and g27077 ( n23159 , n17308 , n31773 );
    not g27078 ( n3191 , n9424 );
    xnor g27079 ( n5570 , n30333 , n23901 );
    or g27080 ( n9004 , n30647 , n2664 );
    and g27081 ( n1801 , n29823 , n85 );
    nor g27082 ( n9290 , n8278 , n28273 );
    or g27083 ( n27463 , n1768 , n22986 );
    not g27084 ( n3021 , n22640 );
    and g27085 ( n24484 , n21887 , n6385 );
    xnor g27086 ( n31336 , n25208 , n18253 );
    not g27087 ( n7764 , n16002 );
    not g27088 ( n1154 , n26956 );
    not g27089 ( n24814 , n27196 );
    not g27090 ( n24548 , n17634 );
    xnor g27091 ( n18914 , n29843 , n6071 );
    not g27092 ( n137 , n27143 );
    nor g27093 ( n24545 , n9375 , n24832 );
    xor g27094 ( n14394 , n883 , n4878 );
    or g27095 ( n113 , n10713 , n9551 );
    not g27096 ( n1461 , n12383 );
    and g27097 ( n4366 , n22362 , n17587 );
    or g27098 ( n2223 , n2989 , n18757 );
    or g27099 ( n26857 , n27052 , n11038 );
    or g27100 ( n1916 , n22406 , n31087 );
    not g27101 ( n10826 , n29441 );
    and g27102 ( n26827 , n24658 , n29019 );
    and g27103 ( n15234 , n1727 , n21172 );
    not g27104 ( n22996 , n10938 );
    or g27105 ( n17874 , n9808 , n28554 );
    not g27106 ( n10081 , n5268 );
    xnor g27107 ( n30541 , n13477 , n10565 );
    or g27108 ( n10247 , n18412 , n5924 );
    xnor g27109 ( n6544 , n14586 , n15715 );
    xnor g27110 ( n22586 , n29257 , n31904 );
    xnor g27111 ( n28903 , n5870 , n736 );
    and g27112 ( n10656 , n28635 , n19211 );
    not g27113 ( n30991 , n10244 );
    not g27114 ( n7457 , n27034 );
    and g27115 ( n24931 , n20580 , n29530 );
    or g27116 ( n29410 , n9204 , n23141 );
    not g27117 ( n18992 , n20980 );
    xnor g27118 ( n4367 , n466 , n14670 );
    xnor g27119 ( n4587 , n29539 , n16061 );
    nor g27120 ( n4824 , n25878 , n23857 );
    and g27121 ( n10307 , n422 , n19903 );
    xnor g27122 ( n3048 , n31316 , n21014 );
    not g27123 ( n19708 , n1205 );
    and g27124 ( n20117 , n11748 , n24883 );
    or g27125 ( n10359 , n16012 , n30809 );
    and g27126 ( n5939 , n14362 , n9338 );
    not g27127 ( n25988 , n10844 );
    not g27128 ( n10328 , n18857 );
    not g27129 ( n2267 , n25413 );
    and g27130 ( n20576 , n8889 , n1836 );
    not g27131 ( n14595 , n23644 );
    xnor g27132 ( n29514 , n9934 , n11755 );
    not g27133 ( n5180 , n17971 );
    and g27134 ( n19552 , n6570 , n22354 );
    or g27135 ( n2099 , n26396 , n209 );
    or g27136 ( n19992 , n8584 , n16716 );
    not g27137 ( n14087 , n23802 );
    not g27138 ( n5974 , n6890 );
    xnor g27139 ( n18832 , n2795 , n31494 );
    not g27140 ( n7352 , n6686 );
    or g27141 ( n15445 , n3302 , n19623 );
    not g27142 ( n3310 , n18305 );
    not g27143 ( n27429 , n20755 );
    not g27144 ( n30629 , n20382 );
    or g27145 ( n10111 , n14364 , n5871 );
    xnor g27146 ( n2062 , n17149 , n20041 );
    not g27147 ( n24392 , n22718 );
    nor g27148 ( n6967 , n23176 , n8506 );
    xnor g27149 ( n6992 , n22511 , n4729 );
    or g27150 ( n791 , n15176 , n6426 );
    nor g27151 ( n27262 , n7763 , n14585 );
    xnor g27152 ( n7830 , n23271 , n12368 );
    and g27153 ( n12891 , n8571 , n24327 );
    xnor g27154 ( n11539 , n16803 , n10393 );
    or g27155 ( n4585 , n17851 , n18042 );
    nor g27156 ( n12716 , n13813 , n6372 );
    not g27157 ( n8234 , n31748 );
    or g27158 ( n10923 , n4956 , n33 );
    not g27159 ( n1410 , n31216 );
    or g27160 ( n10140 , n3977 , n22683 );
    or g27161 ( n582 , n31200 , n2162 );
    or g27162 ( n9804 , n26138 , n13977 );
    or g27163 ( n27804 , n6532 , n8742 );
    xnor g27164 ( n9628 , n4030 , n13549 );
    xnor g27165 ( n3643 , n4335 , n27002 );
    or g27166 ( n16169 , n18493 , n29562 );
    or g27167 ( n3666 , n31730 , n15963 );
    xnor g27168 ( n11363 , n22370 , n13858 );
    not g27169 ( n7390 , n9163 );
    nor g27170 ( n18319 , n24171 , n21066 );
    and g27171 ( n3776 , n3931 , n20847 );
    nor g27172 ( n13530 , n5825 , n28468 );
    nor g27173 ( n1201 , n17609 , n25674 );
    xnor g27174 ( n26379 , n16387 , n7384 );
    or g27175 ( n436 , n19304 , n29899 );
    not g27176 ( n13752 , n11197 );
    or g27177 ( n17908 , n29599 , n21904 );
    or g27178 ( n26574 , n1621 , n26776 );
    not g27179 ( n6775 , n29974 );
    not g27180 ( n21336 , n19348 );
    or g27181 ( n21705 , n1116 , n13455 );
    not g27182 ( n23647 , n28081 );
    or g27183 ( n10945 , n29861 , n21695 );
    not g27184 ( n17909 , n26185 );
    and g27185 ( n5929 , n26782 , n19249 );
    or g27186 ( n16021 , n31685 , n27446 );
    and g27187 ( n8821 , n11553 , n17891 );
    xnor g27188 ( n3937 , n16303 , n13871 );
    or g27189 ( n7581 , n1856 , n14380 );
    or g27190 ( n9017 , n6104 , n7645 );
    not g27191 ( n18464 , n16803 );
    not g27192 ( n8496 , n4588 );
    not g27193 ( n16800 , n2019 );
    not g27194 ( n10374 , n9696 );
    nor g27195 ( n14553 , n21336 , n23567 );
    or g27196 ( n8129 , n32006 , n3927 );
    and g27197 ( n13002 , n29489 , n4842 );
    or g27198 ( n21351 , n25385 , n19324 );
    not g27199 ( n17784 , n18394 );
    or g27200 ( n19798 , n8292 , n25677 );
    xor g27201 ( n11036 , n26225 , n19938 );
    or g27202 ( n10715 , n27618 , n6834 );
    or g27203 ( n17422 , n20487 , n3797 );
    not g27204 ( n14202 , n1177 );
    xnor g27205 ( n17559 , n8939 , n21653 );
    not g27206 ( n6770 , n22743 );
    or g27207 ( n15931 , n9768 , n14969 );
    xnor g27208 ( n25002 , n17247 , n26971 );
    and g27209 ( n1541 , n14636 , n12055 );
    or g27210 ( n26600 , n20836 , n1591 );
    xnor g27211 ( n20593 , n3178 , n31109 );
    not g27212 ( n26969 , n31465 );
    xnor g27213 ( n32021 , n13216 , n23387 );
    or g27214 ( n9273 , n2639 , n145 );
    not g27215 ( n11118 , n7623 );
    and g27216 ( n24061 , n27067 , n31111 );
    xnor g27217 ( n9944 , n17617 , n11789 );
    not g27218 ( n11102 , n9818 );
    not g27219 ( n29891 , n18165 );
    not g27220 ( n7338 , n12630 );
    or g27221 ( n31459 , n15800 , n29423 );
    or g27222 ( n17043 , n3822 , n7414 );
    not g27223 ( n23247 , n30335 );
    not g27224 ( n13300 , n22905 );
    xnor g27225 ( n29747 , n6289 , n17065 );
    nor g27226 ( n4538 , n16982 , n11100 );
    xnor g27227 ( n25125 , n19255 , n8714 );
    xnor g27228 ( n26262 , n14872 , n13725 );
    xnor g27229 ( n6043 , n21840 , n12020 );
    buf g27230 ( n27481 , n27483 );
    not g27231 ( n18776 , n26212 );
    not g27232 ( n25598 , n25938 );
    or g27233 ( n17309 , n4648 , n10658 );
    and g27234 ( n17795 , n31208 , n5645 );
    xor g27235 ( n10172 , n19579 , n11390 );
    not g27236 ( n10348 , n1786 );
    not g27237 ( n18762 , n2287 );
    xnor g27238 ( n25920 , n10058 , n7215 );
    not g27239 ( n23017 , n10738 );
    xnor g27240 ( n9144 , n29501 , n13815 );
    xnor g27241 ( n29593 , n14394 , n10323 );
    xnor g27242 ( n30089 , n22364 , n1401 );
    not g27243 ( n5679 , n6737 );
    and g27244 ( n6348 , n7984 , n26588 );
    not g27245 ( n21407 , n9508 );
    or g27246 ( n1753 , n27376 , n31596 );
    xnor g27247 ( n17491 , n425 , n28589 );
    not g27248 ( n13759 , n11676 );
    and g27249 ( n5527 , n23059 , n12015 );
    xnor g27250 ( n15983 , n18907 , n1995 );
    xnor g27251 ( n24440 , n18750 , n107 );
    not g27252 ( n2527 , n29896 );
    xnor g27253 ( n19856 , n3385 , n11307 );
    not g27254 ( n9216 , n13768 );
    not g27255 ( n6395 , n8134 );
    or g27256 ( n29694 , n14899 , n13101 );
    or g27257 ( n23782 , n30781 , n5722 );
    and g27258 ( n31244 , n30370 , n3163 );
    xnor g27259 ( n1320 , n7209 , n27591 );
    and g27260 ( n28725 , n3220 , n23011 );
    xnor g27261 ( n12727 , n27099 , n9629 );
    buf g27262 ( n16540 , n2185 );
    not g27263 ( n14867 , n4361 );
    not g27264 ( n8845 , n17477 );
    xnor g27265 ( n3523 , n26450 , n1663 );
    not g27266 ( n24018 , n12384 );
    xnor g27267 ( n26947 , n7202 , n15244 );
    xnor g27268 ( n29341 , n8848 , n8654 );
    nor g27269 ( n19376 , n9221 , n9293 );
    and g27270 ( n17344 , n31820 , n7279 );
    not g27271 ( n7336 , n18833 );
    or g27272 ( n21916 , n12954 , n28246 );
    nor g27273 ( n6713 , n28634 , n11641 );
    or g27274 ( n6420 , n21592 , n18347 );
    and g27275 ( n143 , n28175 , n8816 );
    xnor g27276 ( n17111 , n24269 , n30962 );
    or g27277 ( n7759 , n8575 , n22052 );
    not g27278 ( n16599 , n11583 );
    not g27279 ( n30095 , n12199 );
    or g27280 ( n25696 , n19160 , n24254 );
    or g27281 ( n26263 , n11316 , n17738 );
    or g27282 ( n24072 , n1564 , n26970 );
    not g27283 ( n15750 , n28978 );
    xnor g27284 ( n3000 , n17164 , n25585 );
    xnor g27285 ( n21966 , n9020 , n30606 );
    not g27286 ( n519 , n22904 );
    and g27287 ( n29750 , n8851 , n29931 );
    not g27288 ( n26798 , n9124 );
    or g27289 ( n26107 , n25903 , n7966 );
    nor g27290 ( n11853 , n10476 , n18679 );
    xnor g27291 ( n1528 , n26559 , n20400 );
    not g27292 ( n26833 , n7104 );
    or g27293 ( n14622 , n8990 , n8216 );
    not g27294 ( n9285 , n8758 );
    xnor g27295 ( n24618 , n14227 , n19092 );
    or g27296 ( n15326 , n9002 , n20385 );
    xor g27297 ( n4509 , n26060 , n24525 );
    not g27298 ( n6850 , n7798 );
    or g27299 ( n4291 , n22977 , n26633 );
    or g27300 ( n20244 , n9559 , n20849 );
    or g27301 ( n9992 , n17081 , n25223 );
    and g27302 ( n29535 , n9707 , n6312 );
    or g27303 ( n21456 , n19632 , n8166 );
    buf g27304 ( n13888 , n8775 );
    or g27305 ( n5158 , n30514 , n7777 );
    or g27306 ( n19232 , n23620 , n31104 );
    or g27307 ( n9936 , n1983 , n19021 );
    xnor g27308 ( n141 , n6684 , n8847 );
    and g27309 ( n13675 , n15003 , n21251 );
    xnor g27310 ( n20966 , n25621 , n27952 );
    and g27311 ( n28704 , n14574 , n15914 );
    and g27312 ( n29670 , n17841 , n4749 );
    or g27313 ( n8636 , n11295 , n9025 );
    or g27314 ( n25475 , n11883 , n30766 );
    not g27315 ( n14672 , n1718 );
    or g27316 ( n26291 , n23572 , n13451 );
    or g27317 ( n23049 , n11094 , n9461 );
    or g27318 ( n6019 , n23736 , n13158 );
    and g27319 ( n22505 , n156 , n21289 );
    and g27320 ( n174 , n7448 , n19595 );
    xnor g27321 ( n18993 , n16897 , n30142 );
    xnor g27322 ( n23154 , n28165 , n15887 );
    not g27323 ( n24400 , n12139 );
    xnor g27324 ( n20641 , n11999 , n30987 );
    and g27325 ( n15399 , n13752 , n238 );
    xnor g27326 ( n8109 , n3327 , n690 );
    and g27327 ( n5597 , n3860 , n16585 );
    not g27328 ( n16863 , n27971 );
    and g27329 ( n5512 , n4025 , n9344 );
    not g27330 ( n3303 , n16079 );
    or g27331 ( n3467 , n25786 , n20577 );
    or g27332 ( n14283 , n4528 , n31683 );
    xnor g27333 ( n8822 , n31024 , n17171 );
    not g27334 ( n15154 , n19315 );
    not g27335 ( n26235 , n9591 );
    not g27336 ( n29237 , n1396 );
    xnor g27337 ( n15372 , n29960 , n19003 );
    not g27338 ( n26423 , n1119 );
    not g27339 ( n17118 , n23306 );
    not g27340 ( n16833 , n17620 );
    xnor g27341 ( n10389 , n18006 , n31413 );
    or g27342 ( n4616 , n28193 , n293 );
    or g27343 ( n8840 , n11493 , n24288 );
    and g27344 ( n26289 , n26794 , n20181 );
    not g27345 ( n2849 , n20379 );
    or g27346 ( n12670 , n18876 , n6164 );
    not g27347 ( n7998 , n13111 );
    not g27348 ( n9488 , n18855 );
    and g27349 ( n22276 , n7952 , n11750 );
    or g27350 ( n2961 , n21546 , n9054 );
    xnor g27351 ( n6261 , n404 , n13576 );
    and g27352 ( n26589 , n29208 , n30581 );
    or g27353 ( n1864 , n26203 , n10670 );
    or g27354 ( n12947 , n3726 , n16098 );
    not g27355 ( n3350 , n27403 );
    nor g27356 ( n11231 , n14496 , n21934 );
    and g27357 ( n5469 , n13625 , n24163 );
    or g27358 ( n15660 , n6301 , n5694 );
    xnor g27359 ( n12262 , n2543 , n4847 );
    not g27360 ( n28001 , n27764 );
    xnor g27361 ( n19889 , n12192 , n7137 );
    or g27362 ( n12876 , n6534 , n10658 );
    not g27363 ( n25466 , n10323 );
    xnor g27364 ( n298 , n7024 , n12364 );
    or g27365 ( n30843 , n23294 , n7504 );
    and g27366 ( n16194 , n5834 , n3830 );
    or g27367 ( n27078 , n12268 , n29115 );
    and g27368 ( n13384 , n27197 , n19266 );
    xnor g27369 ( n5981 , n14827 , n13952 );
    or g27370 ( n7572 , n31432 , n17300 );
    xnor g27371 ( n8611 , n4786 , n13410 );
    xnor g27372 ( n17832 , n14482 , n6286 );
    nor g27373 ( n23479 , n15667 , n11628 );
    and g27374 ( n425 , n8170 , n2412 );
    not g27375 ( n23652 , n24175 );
    xnor g27376 ( n14665 , n16102 , n24851 );
    and g27377 ( n9955 , n27852 , n24887 );
    and g27378 ( n22239 , n22222 , n15994 );
    xnor g27379 ( n8236 , n14070 , n10955 );
    not g27380 ( n12214 , n1318 );
    or g27381 ( n20287 , n13137 , n20397 );
    not g27382 ( n9279 , n12794 );
    xnor g27383 ( n28154 , n6879 , n9011 );
    and g27384 ( n4180 , n8072 , n30531 );
    xor g27385 ( n4795 , n9021 , n28789 );
    xnor g27386 ( n48 , n14014 , n6952 );
    or g27387 ( n17724 , n19946 , n25241 );
    or g27388 ( n17303 , n13853 , n20523 );
    or g27389 ( n16262 , n28219 , n31155 );
    not g27390 ( n28735 , n24352 );
    not g27391 ( n11198 , n9550 );
    and g27392 ( n14472 , n24108 , n6663 );
    xnor g27393 ( n22087 , n25823 , n9157 );
    xnor g27394 ( n12327 , n10269 , n17255 );
    and g27395 ( n31410 , n6201 , n15938 );
    not g27396 ( n24844 , n8572 );
    nor g27397 ( n15411 , n26750 , n18762 );
    and g27398 ( n19355 , n25826 , n9505 );
    xnor g27399 ( n317 , n4467 , n15822 );
    not g27400 ( n1054 , n31968 );
    or g27401 ( n14596 , n29974 , n5441 );
    not g27402 ( n24049 , n13558 );
    xnor g27403 ( n9585 , n7489 , n5113 );
    not g27404 ( n31953 , n17548 );
    xnor g27405 ( n11949 , n3521 , n22135 );
    or g27406 ( n3474 , n31822 , n10978 );
    xnor g27407 ( n8475 , n21037 , n29580 );
    not g27408 ( n21025 , n26511 );
    xnor g27409 ( n12695 , n19688 , n17492 );
    not g27410 ( n17477 , n13585 );
    and g27411 ( n2823 , n19480 , n25292 );
    xnor g27412 ( n17896 , n31307 , n4393 );
    or g27413 ( n19139 , n20462 , n6408 );
    not g27414 ( n7347 , n181 );
    not g27415 ( n16181 , n23474 );
    and g27416 ( n9126 , n19423 , n22310 );
    xnor g27417 ( n9105 , n6746 , n13876 );
    and g27418 ( n9447 , n19350 , n29025 );
    not g27419 ( n25730 , n16943 );
    nor g27420 ( n21169 , n11132 , n939 );
    xor g27421 ( n26814 , n31835 , n19830 );
    or g27422 ( n10878 , n22144 , n17031 );
    xnor g27423 ( n16830 , n1887 , n6320 );
    not g27424 ( n21158 , n13331 );
    or g27425 ( n22488 , n17098 , n7686 );
    or g27426 ( n23975 , n11601 , n25550 );
    not g27427 ( n16887 , n10404 );
    not g27428 ( n32001 , n27996 );
    or g27429 ( n31442 , n15527 , n28090 );
    and g27430 ( n31054 , n17944 , n28970 );
    or g27431 ( n11529 , n22274 , n17552 );
    or g27432 ( n31932 , n10293 , n30223 );
    not g27433 ( n26843 , n2405 );
    xnor g27434 ( n19671 , n18961 , n20843 );
    xnor g27435 ( n10677 , n23651 , n7180 );
    xnor g27436 ( n21931 , n19005 , n22464 );
    not g27437 ( n1262 , n14021 );
    xnor g27438 ( n16924 , n30505 , n11771 );
    nor g27439 ( n23543 , n867 , n3714 );
    nor g27440 ( n18974 , n15441 , n8801 );
    not g27441 ( n26890 , n14267 );
    xnor g27442 ( n5024 , n13302 , n9673 );
    not g27443 ( n20459 , n29285 );
    or g27444 ( n21051 , n3318 , n23332 );
    nor g27445 ( n5653 , n26365 , n5062 );
    nor g27446 ( n3640 , n10081 , n3267 );
    and g27447 ( n3458 , n17299 , n20278 );
    xnor g27448 ( n4271 , n4312 , n25620 );
    xnor g27449 ( n28272 , n24230 , n11118 );
    not g27450 ( n12596 , n2516 );
    or g27451 ( n29626 , n15589 , n4701 );
    xnor g27452 ( n1309 , n25076 , n8981 );
    not g27453 ( n10069 , n11250 );
    and g27454 ( n14625 , n11382 , n9795 );
    or g27455 ( n31377 , n8912 , n24760 );
    and g27456 ( n16137 , n6450 , n30048 );
    xnor g27457 ( n27571 , n15443 , n9406 );
    or g27458 ( n9953 , n18599 , n10492 );
    and g27459 ( n1749 , n21020 , n30769 );
    xnor g27460 ( n2075 , n31727 , n7354 );
    xnor g27461 ( n22341 , n14992 , n11197 );
    xnor g27462 ( n13760 , n23292 , n7465 );
    or g27463 ( n9314 , n12013 , n24270 );
    or g27464 ( n27933 , n16739 , n6831 );
    xor g27465 ( n7204 , n7777 , n17347 );
    and g27466 ( n14130 , n16606 , n18859 );
    and g27467 ( n24532 , n21566 , n4031 );
    or g27468 ( n10963 , n230 , n23878 );
    not g27469 ( n11468 , n29391 );
    nor g27470 ( n25868 , n12607 , n9987 );
    not g27471 ( n31972 , n26353 );
    not g27472 ( n18143 , n8087 );
    xnor g27473 ( n3935 , n29531 , n24134 );
    not g27474 ( n29226 , n4194 );
    xnor g27475 ( n10407 , n5029 , n29474 );
    not g27476 ( n12080 , n22254 );
    or g27477 ( n13921 , n26419 , n14744 );
    not g27478 ( n19200 , n25335 );
    or g27479 ( n10410 , n7046 , n14266 );
    not g27480 ( n19182 , n6342 );
    xnor g27481 ( n31519 , n28596 , n13205 );
    xnor g27482 ( n1268 , n20229 , n23752 );
    or g27483 ( n30605 , n6189 , n14564 );
    not g27484 ( n23521 , n31882 );
    or g27485 ( n10808 , n19693 , n8577 );
    and g27486 ( n17360 , n21645 , n26994 );
    or g27487 ( n26935 , n19285 , n29267 );
    and g27488 ( n6035 , n18340 , n11083 );
    or g27489 ( n14512 , n4060 , n22458 );
    or g27490 ( n18305 , n6256 , n3435 );
    or g27491 ( n14654 , n31244 , n1907 );
    or g27492 ( n4015 , n11520 , n12371 );
    and g27493 ( n24207 , n24168 , n18923 );
    xnor g27494 ( n31143 , n25 , n17457 );
    or g27495 ( n19501 , n26052 , n4511 );
    xnor g27496 ( n2331 , n6077 , n23041 );
    and g27497 ( n21912 , n27827 , n10954 );
    and g27498 ( n18918 , n16089 , n5222 );
    xnor g27499 ( n3995 , n31065 , n18019 );
    or g27500 ( n26460 , n11662 , n2048 );
    nor g27501 ( n22532 , n29112 , n27216 );
    xnor g27502 ( n19432 , n23805 , n2397 );
    not g27503 ( n3978 , n22235 );
    and g27504 ( n28466 , n19007 , n11226 );
    not g27505 ( n15631 , n20315 );
    xnor g27506 ( n15971 , n10298 , n23571 );
    or g27507 ( n11090 , n23966 , n10899 );
    xnor g27508 ( n20391 , n12242 , n9509 );
    xnor g27509 ( n27085 , n3927 , n22921 );
    not g27510 ( n18121 , n15002 );
    and g27511 ( n19479 , n2900 , n3384 );
    xnor g27512 ( n21311 , n22084 , n4013 );
    and g27513 ( n31392 , n12549 , n20614 );
    xnor g27514 ( n28168 , n21274 , n28569 );
    xnor g27515 ( n13653 , n13091 , n30363 );
    nor g27516 ( n16648 , n10559 , n13723 );
    and g27517 ( n26913 , n18845 , n23221 );
    and g27518 ( n32003 , n1683 , n7131 );
    not g27519 ( n7129 , n11668 );
    xnor g27520 ( n9073 , n20315 , n17210 );
    xnor g27521 ( n12199 , n17709 , n28520 );
    and g27522 ( n26967 , n27712 , n21255 );
    or g27523 ( n21519 , n30688 , n1270 );
    not g27524 ( n3716 , n17531 );
    nor g27525 ( n16592 , n3312 , n21522 );
    or g27526 ( n21593 , n4264 , n12190 );
    nor g27527 ( n248 , n9310 , n4924 );
    not g27528 ( n12740 , n16973 );
    or g27529 ( n882 , n20895 , n4715 );
    or g27530 ( n13078 , n23855 , n16979 );
    nor g27531 ( n31406 , n16779 , n31450 );
    and g27532 ( n14723 , n11426 , n11497 );
    not g27533 ( n16147 , n12143 );
    not g27534 ( n8619 , n29386 );
    and g27535 ( n19297 , n9666 , n7975 );
    not g27536 ( n17295 , n16008 );
    nor g27537 ( n30348 , n13158 , n29867 );
    not g27538 ( n31761 , n14422 );
    or g27539 ( n24556 , n9546 , n9946 );
    not g27540 ( n7182 , n26863 );
    nor g27541 ( n28985 , n8260 , n16637 );
    or g27542 ( n9552 , n21457 , n16797 );
    and g27543 ( n15106 , n5943 , n24872 );
    not g27544 ( n3565 , n24975 );
    xnor g27545 ( n25641 , n5399 , n29972 );
    xnor g27546 ( n23170 , n14672 , n3546 );
    or g27547 ( n27124 , n6613 , n24947 );
    not g27548 ( n17890 , n25076 );
    or g27549 ( n11260 , n12605 , n13486 );
    and g27550 ( n16433 , n10126 , n8373 );
    and g27551 ( n25303 , n23657 , n16084 );
    and g27552 ( n19605 , n16447 , n24395 );
    not g27553 ( n29926 , n11127 );
    xnor g27554 ( n31198 , n24111 , n10841 );
    or g27555 ( n27671 , n8147 , n702 );
    xor g27556 ( n23143 , n540 , n17697 );
    xnor g27557 ( n25553 , n28593 , n28956 );
    xnor g27558 ( n13262 , n25456 , n11719 );
    or g27559 ( n13715 , n17460 , n15798 );
    xnor g27560 ( n8319 , n15404 , n13309 );
    not g27561 ( n13129 , n31988 );
    or g27562 ( n6201 , n24576 , n12267 );
    not g27563 ( n163 , n17184 );
    or g27564 ( n14156 , n28330 , n30841 );
    and g27565 ( n13863 , n12731 , n27051 );
    not g27566 ( n19140 , n27295 );
    or g27567 ( n12769 , n11866 , n551 );
    xnor g27568 ( n6080 , n5587 , n21605 );
    nor g27569 ( n24038 , n13957 , n15819 );
    and g27570 ( n5162 , n27983 , n4746 );
    xnor g27571 ( n17992 , n27644 , n27657 );
    not g27572 ( n2228 , n15448 );
    not g27573 ( n11413 , n15472 );
    and g27574 ( n7591 , n27928 , n20249 );
    or g27575 ( n27561 , n19601 , n26350 );
    or g27576 ( n18695 , n4877 , n28206 );
    nor g27577 ( n662 , n23513 , n13322 );
    or g27578 ( n1959 , n157 , n12719 );
    or g27579 ( n7863 , n6789 , n25680 );
    or g27580 ( n29518 , n27287 , n13636 );
    or g27581 ( n30226 , n31009 , n18780 );
    nor g27582 ( n10554 , n30321 , n16692 );
    not g27583 ( n26161 , n23320 );
    not g27584 ( n25756 , n18416 );
    not g27585 ( n18097 , n2517 );
    not g27586 ( n1730 , n16920 );
    nor g27587 ( n12269 , n20834 , n15262 );
    or g27588 ( n25317 , n29907 , n23629 );
    not g27589 ( n6129 , n25415 );
    or g27590 ( n28163 , n20526 , n13118 );
    xnor g27591 ( n12669 , n23329 , n15538 );
    xnor g27592 ( n28257 , n18486 , n27752 );
    not g27593 ( n1526 , n28460 );
    not g27594 ( n319 , n28614 );
    or g27595 ( n16519 , n18457 , n27024 );
    xnor g27596 ( n16536 , n17 , n13986 );
    xnor g27597 ( n28663 , n8881 , n4218 );
    and g27598 ( n22983 , n1750 , n19501 );
    and g27599 ( n11476 , n16432 , n17193 );
    not g27600 ( n202 , n29323 );
    not g27601 ( n1870 , n9443 );
    not g27602 ( n31880 , n16965 );
    or g27603 ( n19141 , n11360 , n1860 );
    xnor g27604 ( n25601 , n2796 , n1944 );
    not g27605 ( n20299 , n6491 );
    and g27606 ( n6484 , n22162 , n27349 );
    or g27607 ( n4333 , n29332 , n2597 );
    xor g27608 ( n8281 , n7051 , n9096 );
    and g27609 ( n7610 , n24720 , n1357 );
    and g27610 ( n23827 , n11496 , n8353 );
    nor g27611 ( n495 , n10934 , n21307 );
    or g27612 ( n24726 , n17218 , n17086 );
    and g27613 ( n28348 , n1326 , n8016 );
    not g27614 ( n27513 , n20546 );
    not g27615 ( n3530 , n10875 );
    xnor g27616 ( n13457 , n26 , n13249 );
    xnor g27617 ( n30819 , n24939 , n14035 );
    nor g27618 ( n9453 , n14931 , n16867 );
    and g27619 ( n28935 , n28569 , n27473 );
    xnor g27620 ( n28779 , n13918 , n10477 );
    and g27621 ( n6958 , n13069 , n24506 );
    and g27622 ( n10770 , n7490 , n25865 );
    not g27623 ( n9871 , n27733 );
    or g27624 ( n743 , n20049 , n6091 );
    or g27625 ( n23537 , n21969 , n11146 );
    not g27626 ( n11901 , n26846 );
    or g27627 ( n1029 , n2340 , n12741 );
    not g27628 ( n25504 , n31966 );
    or g27629 ( n1596 , n9714 , n18643 );
    xnor g27630 ( n16214 , n7531 , n25746 );
    and g27631 ( n30620 , n29781 , n876 );
    or g27632 ( n22362 , n30193 , n28723 );
    or g27633 ( n24078 , n2009 , n2579 );
    or g27634 ( n9313 , n24334 , n3330 );
    not g27635 ( n29788 , n27692 );
    nor g27636 ( n17570 , n16728 , n11159 );
    not g27637 ( n23092 , n20467 );
    nor g27638 ( n26797 , n1635 , n17330 );
    xnor g27639 ( n21080 , n5063 , n26653 );
    xnor g27640 ( n12597 , n31125 , n30769 );
    or g27641 ( n21575 , n26332 , n1260 );
    or g27642 ( n7888 , n18568 , n910 );
    or g27643 ( n18786 , n1899 , n816 );
    or g27644 ( n17264 , n15681 , n31673 );
    xnor g27645 ( n16500 , n22183 , n1577 );
    xnor g27646 ( n12329 , n12472 , n15417 );
    not g27647 ( n12346 , n13112 );
    or g27648 ( n12819 , n7465 , n5588 );
    not g27649 ( n23117 , n3837 );
    not g27650 ( n8007 , n17756 );
    not g27651 ( n18118 , n10897 );
    xor g27652 ( n1377 , n21946 , n31818 );
    nor g27653 ( n31234 , n26786 , n1526 );
    or g27654 ( n24603 , n5814 , n16674 );
    not g27655 ( n26569 , n15803 );
    not g27656 ( n30786 , n18943 );
    nor g27657 ( n5804 , n25996 , n21011 );
    or g27658 ( n3165 , n23379 , n30345 );
    nor g27659 ( n30684 , n21275 , n820 );
    not g27660 ( n11047 , n14955 );
    not g27661 ( n21875 , n28815 );
    not g27662 ( n5098 , n2991 );
    or g27663 ( n12484 , n26342 , n3878 );
    and g27664 ( n29329 , n4905 , n27393 );
    xnor g27665 ( n24443 , n20962 , n5073 );
    xnor g27666 ( n19496 , n15554 , n20909 );
    or g27667 ( n30225 , n28365 , n16593 );
    not g27668 ( n10681 , n9176 );
    or g27669 ( n12235 , n6405 , n1446 );
    and g27670 ( n7012 , n10633 , n2447 );
    or g27671 ( n23619 , n2164 , n20398 );
    and g27672 ( n5355 , n31188 , n29615 );
    or g27673 ( n3321 , n24539 , n20742 );
    nor g27674 ( n22619 , n25425 , n16330 );
    or g27675 ( n24240 , n25427 , n31846 );
    not g27676 ( n11745 , n7818 );
    xnor g27677 ( n3888 , n19423 , n28160 );
    not g27678 ( n28407 , n11507 );
    or g27679 ( n10621 , n23320 , n24289 );
    not g27680 ( n4253 , n30586 );
    xnor g27681 ( n11685 , n18656 , n973 );
    xnor g27682 ( n6768 , n22045 , n18380 );
    not g27683 ( n6279 , n9901 );
    xnor g27684 ( n2840 , n1649 , n22184 );
    or g27685 ( n11086 , n24728 , n10355 );
    and g27686 ( n2052 , n3608 , n14541 );
    xnor g27687 ( n6111 , n4359 , n12035 );
    and g27688 ( n10175 , n25722 , n6624 );
    or g27689 ( n23841 , n13638 , n5929 );
    not g27690 ( n26454 , n26758 );
    and g27691 ( n1772 , n12270 , n16515 );
    or g27692 ( n884 , n26777 , n2143 );
    and g27693 ( n4283 , n570 , n26730 );
    xnor g27694 ( n31477 , n2890 , n11445 );
    not g27695 ( n2689 , n12980 );
    not g27696 ( n8865 , n1120 );
    nor g27697 ( n30515 , n22255 , n3558 );
    nor g27698 ( n21395 , n3106 , n14432 );
    xnor g27699 ( n27529 , n2250 , n30391 );
    or g27700 ( n3220 , n9453 , n28171 );
    not g27701 ( n1993 , n27233 );
    not g27702 ( n10367 , n31951 );
    or g27703 ( n1330 , n23576 , n15898 );
    nor g27704 ( n21899 , n27470 , n22382 );
    or g27705 ( n11588 , n10831 , n19872 );
    xnor g27706 ( n599 , n11452 , n27233 );
    not g27707 ( n7143 , n25023 );
    not g27708 ( n21119 , n31546 );
    nor g27709 ( n23162 , n29475 , n31728 );
    xnor g27710 ( n11973 , n18425 , n3688 );
    not g27711 ( n6018 , n32010 );
    nor g27712 ( n3909 , n1935 , n23681 );
    not g27713 ( n31218 , n8238 );
    not g27714 ( n31752 , n29879 );
    not g27715 ( n29131 , n26284 );
    nor g27716 ( n16183 , n23960 , n8586 );
    not g27717 ( n6460 , n17491 );
    or g27718 ( n26111 , n25668 , n31414 );
    not g27719 ( n27965 , n15178 );
    xnor g27720 ( n26065 , n7241 , n19572 );
    not g27721 ( n15145 , n804 );
    nor g27722 ( n18809 , n5675 , n5345 );
    or g27723 ( n30571 , n22382 , n9187 );
    nor g27724 ( n6516 , n24578 , n20390 );
    nor g27725 ( n10290 , n31019 , n7760 );
    not g27726 ( n19383 , n18852 );
    not g27727 ( n479 , n27786 );
    nor g27728 ( n5189 , n20495 , n30088 );
    not g27729 ( n3047 , n28749 );
    and g27730 ( n23166 , n3819 , n13608 );
    not g27731 ( n22977 , n13700 );
    or g27732 ( n22644 , n12889 , n19730 );
    not g27733 ( n17612 , n8934 );
    or g27734 ( n1003 , n8796 , n25087 );
    or g27735 ( n19413 , n6735 , n16845 );
    or g27736 ( n19972 , n30516 , n6043 );
    xnor g27737 ( n21453 , n28246 , n1837 );
    or g27738 ( n20317 , n23195 , n25776 );
    and g27739 ( n15469 , n3685 , n4156 );
    xor g27740 ( n29349 , n631 , n27181 );
    not g27741 ( n23773 , n1770 );
    xnor g27742 ( n3100 , n18921 , n24352 );
    not g27743 ( n22113 , n31313 );
    or g27744 ( n5094 , n24029 , n14660 );
    not g27745 ( n31424 , n3262 );
    not g27746 ( n17834 , n11596 );
    xnor g27747 ( n25952 , n22561 , n842 );
    and g27748 ( n10205 , n8501 , n14301 );
    xor g27749 ( n752 , n30015 , n24321 );
    and g27750 ( n6973 , n22070 , n4991 );
    xnor g27751 ( n18749 , n11629 , n29839 );
    xnor g27752 ( n23483 , n28433 , n16856 );
    xnor g27753 ( n4593 , n21273 , n9724 );
    not g27754 ( n14475 , n22922 );
    nor g27755 ( n8295 , n26929 , n1704 );
    and g27756 ( n16330 , n2267 , n11117 );
    or g27757 ( n8332 , n28673 , n3215 );
    and g27758 ( n2144 , n8657 , n29132 );
    xnor g27759 ( n16981 , n8071 , n16998 );
    and g27760 ( n24208 , n26405 , n14587 );
    and g27761 ( n5554 , n26015 , n3882 );
    buf g27762 ( n2799 , n7162 );
    not g27763 ( n4398 , n29906 );
    and g27764 ( n19618 , n6844 , n32031 );
    nor g27765 ( n419 , n19880 , n775 );
    not g27766 ( n18724 , n21244 );
    or g27767 ( n8721 , n5563 , n7325 );
    xnor g27768 ( n12814 , n10901 , n32004 );
    xnor g27769 ( n28703 , n15801 , n25895 );
    not g27770 ( n31797 , n8407 );
    not g27771 ( n17558 , n9116 );
    or g27772 ( n13379 , n23023 , n13346 );
    not g27773 ( n2842 , n23115 );
    xor g27774 ( n1760 , n7562 , n22525 );
    and g27775 ( n13848 , n26719 , n3835 );
    not g27776 ( n1915 , n6196 );
    xnor g27777 ( n22456 , n3814 , n12305 );
    xnor g27778 ( n29399 , n22366 , n6696 );
    xnor g27779 ( n14883 , n19684 , n18803 );
    and g27780 ( n30947 , n17455 , n12514 );
    and g27781 ( n6373 , n8933 , n3145 );
    not g27782 ( n26647 , n5514 );
    not g27783 ( n20858 , n24299 );
    xnor g27784 ( n30735 , n13865 , n13267 );
    and g27785 ( n17381 , n6460 , n3077 );
    nor g27786 ( n15182 , n22646 , n10759 );
    and g27787 ( n8984 , n22990 , n21593 );
    nor g27788 ( n24966 , n29291 , n31044 );
    or g27789 ( n7074 , n21333 , n14790 );
    or g27790 ( n2039 , n11815 , n4579 );
    nor g27791 ( n19637 , n5149 , n10185 );
    not g27792 ( n28185 , n949 );
    or g27793 ( n8759 , n13753 , n30520 );
    xnor g27794 ( n2024 , n20131 , n31783 );
    or g27795 ( n898 , n8149 , n21944 );
    or g27796 ( n12635 , n19101 , n21137 );
    and g27797 ( n25777 , n14512 , n25816 );
    or g27798 ( n21738 , n30562 , n29118 );
    xnor g27799 ( n23739 , n6395 , n18763 );
    not g27800 ( n4484 , n30916 );
    and g27801 ( n26016 , n342 , n11134 );
    xnor g27802 ( n2170 , n15070 , n1361 );
    not g27803 ( n7385 , n16873 );
    not g27804 ( n23205 , n25026 );
    or g27805 ( n4512 , n8042 , n24527 );
    not g27806 ( n2060 , n19443 );
    or g27807 ( n2790 , n12333 , n19721 );
    or g27808 ( n16577 , n2755 , n7744 );
    not g27809 ( n13132 , n21831 );
    not g27810 ( n22306 , n18763 );
    not g27811 ( n31260 , n1588 );
    nor g27812 ( n10343 , n30931 , n31732 );
    or g27813 ( n7937 , n12837 , n3862 );
    xnor g27814 ( n2691 , n7979 , n29660 );
    and g27815 ( n9601 , n25923 , n28488 );
    xnor g27816 ( n8318 , n11966 , n19755 );
    and g27817 ( n27495 , n9247 , n21065 );
    or g27818 ( n30452 , n7175 , n14833 );
    or g27819 ( n4103 , n21466 , n17995 );
    or g27820 ( n23924 , n31140 , n2723 );
    xnor g27821 ( n6838 , n9414 , n10981 );
    or g27822 ( n27032 , n26236 , n16695 );
    and g27823 ( n23781 , n24316 , n15702 );
    not g27824 ( n8578 , n16602 );
    xnor g27825 ( n2459 , n16838 , n21467 );
    nor g27826 ( n17791 , n6370 , n19777 );
    xnor g27827 ( n15943 , n23471 , n14491 );
    or g27828 ( n15188 , n13279 , n19240 );
    nor g27829 ( n26021 , n22332 , n23335 );
    and g27830 ( n3409 , n8843 , n15601 );
    nor g27831 ( n3242 , n4662 , n5471 );
    or g27832 ( n18600 , n1561 , n10988 );
    not g27833 ( n27690 , n16068 );
    not g27834 ( n10788 , n28035 );
    and g27835 ( n28565 , n15283 , n18302 );
    not g27836 ( n19820 , n7655 );
    and g27837 ( n26968 , n18936 , n29355 );
    xnor g27838 ( n22305 , n20099 , n26231 );
    or g27839 ( n18314 , n10619 , n14324 );
    and g27840 ( n6485 , n19800 , n22327 );
    nor g27841 ( n23674 , n13888 , n2067 );
    or g27842 ( n3334 , n5059 , n17113 );
    xor g27843 ( n8338 , n25229 , n20296 );
    and g27844 ( n13269 , n19463 , n28407 );
    not g27845 ( n25426 , n22330 );
    or g27846 ( n1584 , n20876 , n6242 );
    and g27847 ( n26514 , n29794 , n575 );
    and g27848 ( n29503 , n23468 , n19913 );
    not g27849 ( n17525 , n887 );
    or g27850 ( n22837 , n18941 , n29287 );
    and g27851 ( n27703 , n26480 , n11055 );
    not g27852 ( n14427 , n12783 );
    not g27853 ( n16607 , n7187 );
    not g27854 ( n16404 , n12692 );
    or g27855 ( n19438 , n28351 , n26221 );
    or g27856 ( n7016 , n8834 , n4817 );
    and g27857 ( n14833 , n23384 , n1599 );
    or g27858 ( n7061 , n28172 , n15280 );
    or g27859 ( n11553 , n16866 , n7805 );
    xor g27860 ( n12273 , n997 , n23284 );
    or g27861 ( n9096 , n3828 , n14504 );
    not g27862 ( n4513 , n29647 );
    not g27863 ( n13676 , n26033 );
    nor g27864 ( n28482 , n25031 , n14083 );
    xor g27865 ( n22358 , n4320 , n14611 );
    not g27866 ( n23372 , n17460 );
    not g27867 ( n14538 , n275 );
    or g27868 ( n3551 , n8274 , n25183 );
    and g27869 ( n31387 , n14198 , n27591 );
    not g27870 ( n26351 , n23360 );
    and g27871 ( n10616 , n26276 , n2789 );
    not g27872 ( n14544 , n13502 );
    not g27873 ( n17059 , n31916 );
    nor g27874 ( n9768 , n6141 , n6872 );
    xor g27875 ( n4168 , n2875 , n17137 );
    xnor g27876 ( n13870 , n21394 , n17302 );
    or g27877 ( n7627 , n26089 , n19660 );
    xor g27878 ( n20883 , n8247 , n29480 );
    xnor g27879 ( n7564 , n18492 , n2642 );
    xnor g27880 ( n14712 , n20100 , n12826 );
    and g27881 ( n23065 , n22328 , n1462 );
    not g27882 ( n4075 , n7638 );
    or g27883 ( n22926 , n12276 , n23078 );
    or g27884 ( n11395 , n28731 , n25287 );
    not g27885 ( n22415 , n3303 );
    and g27886 ( n12633 , n17022 , n22672 );
    xnor g27887 ( n18726 , n21007 , n2704 );
    not g27888 ( n8649 , n16890 );
    xnor g27889 ( n14926 , n2225 , n2825 );
    or g27890 ( n31941 , n29400 , n1977 );
    or g27891 ( n5321 , n5313 , n20639 );
    not g27892 ( n31270 , n16536 );
    not g27893 ( n21221 , n15262 );
    nor g27894 ( n5033 , n11974 , n2216 );
    not g27895 ( n21154 , n2128 );
    or g27896 ( n17679 , n8321 , n21442 );
    xnor g27897 ( n19397 , n18926 , n9145 );
    or g27898 ( n17388 , n12290 , n7913 );
    xnor g27899 ( n18685 , n7925 , n16540 );
    not g27900 ( n21667 , n28983 );
    or g27901 ( n28816 , n10840 , n6506 );
    and g27902 ( n24257 , n22815 , n28300 );
    xnor g27903 ( n28237 , n16753 , n12535 );
    not g27904 ( n24913 , n7781 );
    or g27905 ( n4867 , n15645 , n14897 );
    and g27906 ( n9504 , n17984 , n13715 );
    not g27907 ( n23471 , n24305 );
    nor g27908 ( n18142 , n30664 , n22301 );
    nor g27909 ( n17934 , n8807 , n4695 );
    not g27910 ( n14114 , n29649 );
    and g27911 ( n18828 , n11383 , n21426 );
    xnor g27912 ( n5085 , n28555 , n12832 );
    xnor g27913 ( n15510 , n83 , n15946 );
    xnor g27914 ( n19965 , n4462 , n25618 );
    nor g27915 ( n3149 , n1845 , n29326 );
    and g27916 ( n28157 , n29819 , n11384 );
    or g27917 ( n27912 , n13766 , n19834 );
    not g27918 ( n23271 , n5818 );
    not g27919 ( n29663 , n24540 );
    nor g27920 ( n18239 , n30254 , n10068 );
    xnor g27921 ( n11752 , n3765 , n14992 );
    nor g27922 ( n28329 , n11101 , n9718 );
    or g27923 ( n4792 , n16771 , n16257 );
    and g27924 ( n3766 , n13873 , n23981 );
    not g27925 ( n12772 , n28384 );
    xnor g27926 ( n23486 , n29825 , n15552 );
    not g27927 ( n10710 , n14233 );
    and g27928 ( n31876 , n31093 , n23386 );
    nor g27929 ( n15888 , n7781 , n24322 );
    xnor g27930 ( n12790 , n25354 , n25337 );
    and g27931 ( n27623 , n2707 , n9977 );
    nor g27932 ( n21344 , n1616 , n21597 );
    nor g27933 ( n4147 , n1935 , n16238 );
    not g27934 ( n14480 , n23738 );
    xnor g27935 ( n28860 , n5608 , n8483 );
    or g27936 ( n31216 , n28280 , n20109 );
    or g27937 ( n11978 , n2894 , n3067 );
    xnor g27938 ( n24980 , n10114 , n3782 );
    and g27939 ( n9191 , n13742 , n6344 );
    and g27940 ( n838 , n10337 , n23515 );
    not g27941 ( n5788 , n4554 );
    and g27942 ( n28078 , n24308 , n5570 );
    xnor g27943 ( n5455 , n19451 , n2313 );
    not g27944 ( n10533 , n25629 );
    not g27945 ( n25045 , n26058 );
    nor g27946 ( n14420 , n22631 , n30131 );
    not g27947 ( n11983 , n15550 );
    not g27948 ( n23002 , n28121 );
    not g27949 ( n12428 , n6957 );
    or g27950 ( n7166 , n19632 , n26852 );
    not g27951 ( n29591 , n10042 );
    not g27952 ( n19597 , n29248 );
    not g27953 ( n27012 , n7021 );
    not g27954 ( n18045 , n7009 );
    and g27955 ( n12534 , n9992 , n3049 );
    nor g27956 ( n2705 , n16338 , n24405 );
    or g27957 ( n2455 , n22910 , n28430 );
    not g27958 ( n23628 , n27521 );
    or g27959 ( n16961 , n14711 , n25827 );
    or g27960 ( n9331 , n15367 , n27634 );
    xnor g27961 ( n26470 , n18186 , n21533 );
    or g27962 ( n1852 , n21196 , n11196 );
    not g27963 ( n20921 , n8896 );
    not g27964 ( n15737 , n7381 );
    or g27965 ( n22880 , n23639 , n1507 );
    nor g27966 ( n26808 , n31866 , n29366 );
    nor g27967 ( n18377 , n27481 , n14372 );
    xnor g27968 ( n20114 , n11954 , n15147 );
    not g27969 ( n2227 , n27974 );
    and g27970 ( n22770 , n4112 , n16798 );
    not g27971 ( n12493 , n6866 );
    or g27972 ( n5602 , n13372 , n23129 );
    nor g27973 ( n4119 , n28741 , n14825 );
    xnor g27974 ( n13359 , n6656 , n10706 );
    not g27975 ( n6276 , n19857 );
    xnor g27976 ( n22443 , n11680 , n5926 );
    nor g27977 ( n531 , n8018 , n11704 );
    not g27978 ( n25887 , n28666 );
    or g27979 ( n3835 , n13552 , n31372 );
    not g27980 ( n19803 , n10363 );
    not g27981 ( n21059 , n14005 );
    or g27982 ( n22280 , n18239 , n11489 );
    xnor g27983 ( n23414 , n25346 , n18452 );
    not g27984 ( n28912 , n29803 );
    xnor g27985 ( n12699 , n4158 , n19852 );
    xnor g27986 ( n29089 , n10752 , n11405 );
    xor g27987 ( n14392 , n11540 , n22614 );
    not g27988 ( n23900 , n30919 );
    xnor g27989 ( n20518 , n20474 , n22922 );
    xnor g27990 ( n29093 , n28501 , n3734 );
    or g27991 ( n10758 , n13725 , n31361 );
    or g27992 ( n31950 , n1441 , n26546 );
    or g27993 ( n13439 , n27654 , n28266 );
    or g27994 ( n29985 , n8081 , n22086 );
    or g27995 ( n24317 , n177 , n31568 );
    not g27996 ( n3758 , n8890 );
    or g27997 ( n28608 , n15328 , n17424 );
    or g27998 ( n2743 , n25209 , n31230 );
    or g27999 ( n325 , n18862 , n18272 );
    not g28000 ( n10519 , n30958 );
    xnor g28001 ( n8426 , n16564 , n21217 );
    nor g28002 ( n19465 , n21122 , n22135 );
    or g28003 ( n2475 , n16884 , n3919 );
    and g28004 ( n29270 , n8347 , n15762 );
    and g28005 ( n30407 , n3499 , n1986 );
    xor g28006 ( n1501 , n1349 , n12998 );
    not g28007 ( n27473 , n7575 );
    xnor g28008 ( n19648 , n18554 , n8790 );
    not g28009 ( n7230 , n29042 );
    nor g28010 ( n26031 , n6018 , n11944 );
    or g28011 ( n7361 , n18427 , n22110 );
    or g28012 ( n3699 , n30533 , n19758 );
    xnor g28013 ( n14980 , n10848 , n22381 );
    not g28014 ( n28189 , n17069 );
    xnor g28015 ( n6512 , n22147 , n1314 );
    and g28016 ( n21516 , n24042 , n13778 );
    buf g28017 ( n14100 , n25947 );
    not g28018 ( n14162 , n90 );
    and g28019 ( n11200 , n16756 , n22678 );
    xnor g28020 ( n29387 , n21506 , n6689 );
    nor g28021 ( n29107 , n26377 , n13338 );
    and g28022 ( n21015 , n12067 , n22266 );
    or g28023 ( n30280 , n27829 , n1039 );
    not g28024 ( n3535 , n4505 );
    xnor g28025 ( n20437 , n9285 , n30158 );
    or g28026 ( n7403 , n23641 , n5369 );
    or g28027 ( n5850 , n31773 , n13292 );
    not g28028 ( n16254 , n9350 );
    not g28029 ( n7011 , n28426 );
    and g28030 ( n29453 , n4123 , n26937 );
    or g28031 ( n25205 , n13058 , n30870 );
    or g28032 ( n24604 , n30553 , n27525 );
    xnor g28033 ( n23270 , n5830 , n17023 );
    not g28034 ( n1234 , n1021 );
    nor g28035 ( n15727 , n14356 , n8763 );
    xnor g28036 ( n4418 , n28946 , n5792 );
    not g28037 ( n23964 , n2960 );
    not g28038 ( n1650 , n27804 );
    or g28039 ( n24945 , n14987 , n5506 );
    xnor g28040 ( n30142 , n1176 , n11798 );
    xnor g28041 ( n8654 , n29018 , n18 );
    or g28042 ( n9149 , n9737 , n10205 );
    or g28043 ( n24509 , n3688 , n26235 );
    not g28044 ( n23813 , n9152 );
    or g28045 ( n25963 , n18500 , n1650 );
    and g28046 ( n21090 , n349 , n4705 );
    or g28047 ( n26608 , n3837 , n24086 );
    not g28048 ( n30419 , n18511 );
    xnor g28049 ( n1451 , n10557 , n14324 );
    nor g28050 ( n11347 , n25242 , n30135 );
    or g28051 ( n29459 , n4824 , n8082 );
    not g28052 ( n28736 , n9414 );
    or g28053 ( n29501 , n7065 , n24406 );
    and g28054 ( n26110 , n1395 , n30728 );
    xnor g28055 ( n5271 , n25036 , n24820 );
    xnor g28056 ( n2403 , n23311 , n1283 );
    and g28057 ( n7689 , n12791 , n17064 );
    not g28058 ( n28362 , n24798 );
    and g28059 ( n24406 , n27445 , n16876 );
    and g28060 ( n8891 , n29055 , n24002 );
    xnor g28061 ( n15574 , n26687 , n6696 );
    or g28062 ( n16646 , n15035 , n3593 );
    and g28063 ( n29246 , n22556 , n25836 );
    or g28064 ( n6863 , n14535 , n22749 );
    nor g28065 ( n5056 , n16689 , n9137 );
    nor g28066 ( n18944 , n28041 , n22676 );
    xnor g28067 ( n21355 , n13548 , n18133 );
    not g28068 ( n4695 , n21068 );
    not g28069 ( n30560 , n5193 );
    xnor g28070 ( n16412 , n7222 , n3482 );
    and g28071 ( n21413 , n26172 , n9732 );
    nor g28072 ( n5716 , n8853 , n208 );
    or g28073 ( n10478 , n25146 , n2175 );
    and g28074 ( n16303 , n22988 , n17933 );
    nor g28075 ( n9712 , n7729 , n17180 );
    not g28076 ( n4237 , n9353 );
    not g28077 ( n27539 , n26321 );
    and g28078 ( n23067 , n6662 , n28584 );
    or g28079 ( n28488 , n3297 , n31483 );
    xnor g28080 ( n660 , n28381 , n6097 );
    xnor g28081 ( n7779 , n3848 , n6992 );
    nor g28082 ( n5890 , n2352 , n25233 );
    not g28083 ( n4085 , n2599 );
    not g28084 ( n7542 , n4202 );
    not g28085 ( n1568 , n28907 );
    and g28086 ( n18759 , n17322 , n14795 );
    and g28087 ( n14038 , n31532 , n27815 );
    and g28088 ( n6085 , n3650 , n6363 );
    xor g28089 ( n15252 , n7018 , n18988 );
    xnor g28090 ( n14918 , n5831 , n19720 );
    or g28091 ( n22790 , n5388 , n657 );
    not g28092 ( n5853 , n10394 );
    and g28093 ( n31786 , n14448 , n3434 );
    and g28094 ( n18824 , n26868 , n11318 );
    not g28095 ( n30402 , n28502 );
    not g28096 ( n8187 , n29059 );
    nor g28097 ( n8968 , n22079 , n21305 );
    xnor g28098 ( n14316 , n12987 , n27993 );
    or g28099 ( n18304 , n20626 , n1876 );
    not g28100 ( n6509 , n20148 );
    xnor g28101 ( n3928 , n21953 , n2532 );
    nor g28102 ( n7321 , n22912 , n6758 );
    not g28103 ( n28159 , n9739 );
    xnor g28104 ( n1653 , n11396 , n22590 );
    or g28105 ( n19978 , n19514 , n3107 );
    or g28106 ( n10422 , n31185 , n10848 );
    or g28107 ( n30436 , n13123 , n7397 );
    nor g28108 ( n25077 , n15999 , n28962 );
    xnor g28109 ( n30925 , n13408 , n28719 );
    and g28110 ( n7494 , n17500 , n6741 );
    not g28111 ( n23567 , n5261 );
    and g28112 ( n3413 , n30299 , n31774 );
    or g28113 ( n15353 , n9835 , n15620 );
    or g28114 ( n2355 , n10455 , n8367 );
    and g28115 ( n10076 , n10710 , n2798 );
    or g28116 ( n31742 , n24301 , n24967 );
    or g28117 ( n12250 , n20064 , n14760 );
    not g28118 ( n19046 , n19590 );
    xnor g28119 ( n18071 , n13595 , n19124 );
    xnor g28120 ( n21833 , n31405 , n9369 );
    xnor g28121 ( n28470 , n6530 , n28216 );
    and g28122 ( n502 , n13668 , n20608 );
    xnor g28123 ( n7392 , n664 , n29249 );
    nor g28124 ( n13151 , n25699 , n3639 );
    and g28125 ( n16645 , n31248 , n11262 );
    and g28126 ( n12406 , n26900 , n23054 );
    or g28127 ( n22430 , n19035 , n26266 );
    and g28128 ( n13229 , n7100 , n15740 );
    not g28129 ( n4080 , n26372 );
    not g28130 ( n16198 , n24449 );
    and g28131 ( n28910 , n27887 , n25410 );
    not g28132 ( n16453 , n21480 );
    and g28133 ( n13892 , n10425 , n5333 );
    or g28134 ( n26293 , n15004 , n8288 );
    or g28135 ( n8886 , n855 , n6279 );
    or g28136 ( n21190 , n8377 , n18942 );
    xnor g28137 ( n17094 , n27996 , n10888 );
    not g28138 ( n5683 , n2646 );
    not g28139 ( n8453 , n5075 );
    not g28140 ( n2097 , n20218 );
    not g28141 ( n3218 , n26603 );
    or g28142 ( n9003 , n852 , n23293 );
    nor g28143 ( n13938 , n6117 , n29324 );
    not g28144 ( n30229 , n12440 );
    not g28145 ( n7254 , n9217 );
    xnor g28146 ( n13842 , n23665 , n2987 );
    or g28147 ( n5639 , n23487 , n5415 );
    buf g28148 ( n9146 , n28872 );
    not g28149 ( n12489 , n20390 );
    or g28150 ( n16022 , n22914 , n24968 );
    and g28151 ( n3695 , n10111 , n30168 );
    not g28152 ( n28614 , n19393 );
    xnor g28153 ( n11349 , n29622 , n19883 );
    xor g28154 ( n28799 , n4884 , n17328 );
    xnor g28155 ( n19410 , n25302 , n22412 );
    and g28156 ( n23493 , n21690 , n14792 );
    not g28157 ( n10606 , n11630 );
    and g28158 ( n22795 , n20840 , n22584 );
    and g28159 ( n20090 , n14453 , n31962 );
    xnor g28160 ( n16239 , n7374 , n27772 );
    or g28161 ( n24722 , n25113 , n3097 );
    or g28162 ( n29882 , n16137 , n28335 );
    not g28163 ( n31232 , n11101 );
    not g28164 ( n25789 , n27432 );
    or g28165 ( n9437 , n31885 , n12524 );
    not g28166 ( n26945 , n24577 );
    not g28167 ( n26792 , n8680 );
    nor g28168 ( n2954 , n14035 , n154 );
    not g28169 ( n21373 , n2984 );
    and g28170 ( n15556 , n6392 , n29255 );
    not g28171 ( n2067 , n3069 );
    xnor g28172 ( n15286 , n26767 , n15022 );
    xnor g28173 ( n22064 , n7395 , n10388 );
    not g28174 ( n18442 , n31535 );
    nor g28175 ( n13131 , n31910 , n4658 );
    not g28176 ( n19017 , n22377 );
    and g28177 ( n20454 , n25345 , n19430 );
    or g28178 ( n29032 , n9786 , n7126 );
    or g28179 ( n19483 , n13589 , n2332 );
    xnor g28180 ( n21510 , n18936 , n29355 );
    nor g28181 ( n20059 , n14713 , n28987 );
    not g28182 ( n3256 , n29409 );
    nor g28183 ( n27108 , n344 , n20200 );
    and g28184 ( n11151 , n13569 , n26370 );
    xnor g28185 ( n30329 , n10092 , n7650 );
    xnor g28186 ( n17726 , n11796 , n10485 );
    not g28187 ( n26973 , n12701 );
    not g28188 ( n3151 , n8110 );
    not g28189 ( n4758 , n16535 );
    nor g28190 ( n2226 , n20198 , n27549 );
    not g28191 ( n7290 , n28269 );
    nor g28192 ( n1866 , n26451 , n22326 );
    nor g28193 ( n19168 , n15470 , n21564 );
    nor g28194 ( n20282 , n29132 , n16424 );
    not g28195 ( n12580 , n28535 );
    and g28196 ( n12551 , n4452 , n21127 );
    not g28197 ( n11400 , n28427 );
    nor g28198 ( n31767 , n29395 , n26707 );
    or g28199 ( n18294 , n25023 , n22246 );
    not g28200 ( n4498 , n31389 );
    xnor g28201 ( n1360 , n19132 , n18518 );
    not g28202 ( n28449 , n508 );
    or g28203 ( n65 , n14003 , n28360 );
    nor g28204 ( n12002 , n13935 , n17322 );
    or g28205 ( n1816 , n9430 , n9688 );
    not g28206 ( n30314 , n16683 );
    xnor g28207 ( n4694 , n24095 , n19743 );
    and g28208 ( n4463 , n23958 , n17702 );
    xnor g28209 ( n13406 , n22494 , n17094 );
    not g28210 ( n12747 , n14940 );
    or g28211 ( n27907 , n18330 , n26170 );
    xnor g28212 ( n26055 , n30177 , n97 );
    or g28213 ( n5184 , n16630 , n18160 );
    xnor g28214 ( n26790 , n13145 , n25991 );
    not g28215 ( n9889 , n20759 );
    or g28216 ( n7221 , n3736 , n19954 );
    and g28217 ( n29689 , n26680 , n27620 );
    xnor g28218 ( n20662 , n5338 , n25189 );
    and g28219 ( n27991 , n8138 , n16206 );
    not g28220 ( n6995 , n9163 );
    and g28221 ( n1672 , n2333 , n5300 );
    nor g28222 ( n180 , n28154 , n31211 );
    xnor g28223 ( n9479 , n19139 , n22385 );
    not g28224 ( n3821 , n17000 );
    not g28225 ( n6475 , n15631 );
    and g28226 ( n14600 , n23612 , n23020 );
    not g28227 ( n6084 , n24087 );
    not g28228 ( n6960 , n12856 );
    not g28229 ( n26754 , n23236 );
    or g28230 ( n28187 , n27775 , n30574 );
    xnor g28231 ( n7371 , n1156 , n7179 );
    or g28232 ( n9032 , n22528 , n8577 );
    xnor g28233 ( n18435 , n8070 , n29672 );
    or g28234 ( n24453 , n16581 , n18943 );
    not g28235 ( n13822 , n19505 );
    and g28236 ( n21163 , n7702 , n22616 );
    nor g28237 ( n22555 , n9812 , n24381 );
    nor g28238 ( n16712 , n14624 , n7357 );
    not g28239 ( n26587 , n7851 );
    or g28240 ( n30796 , n5936 , n16774 );
    xnor g28241 ( n28512 , n27060 , n8983 );
    xnor g28242 ( n24131 , n5520 , n8639 );
    xnor g28243 ( n29833 , n29235 , n10724 );
    not g28244 ( n12232 , n30649 );
    or g28245 ( n17395 , n12397 , n15547 );
    xnor g28246 ( n26620 , n16480 , n21614 );
    nor g28247 ( n4527 , n5873 , n7229 );
    or g28248 ( n18523 , n31107 , n10141 );
    xnor g28249 ( n16470 , n16113 , n14106 );
    or g28250 ( n13320 , n11713 , n24806 );
    xnor g28251 ( n29229 , n11606 , n24777 );
    not g28252 ( n21363 , n12481 );
    not g28253 ( n20148 , n15017 );
    or g28254 ( n833 , n1863 , n7867 );
    xnor g28255 ( n15855 , n19829 , n8 );
    not g28256 ( n27971 , n15101 );
    not g28257 ( n25436 , n3404 );
    nor g28258 ( n9464 , n17302 , n24969 );
    and g28259 ( n14256 , n12514 , n26456 );
    or g28260 ( n14047 , n10083 , n22336 );
    not g28261 ( n28742 , n6399 );
    xnor g28262 ( n22871 , n568 , n11729 );
    not g28263 ( n14451 , n20105 );
    xnor g28264 ( n1115 , n29970 , n28464 );
    or g28265 ( n22701 , n237 , n20499 );
    not g28266 ( n7200 , n25343 );
    and g28267 ( n23008 , n31209 , n27499 );
    and g28268 ( n23668 , n26673 , n16902 );
    and g28269 ( n21112 , n9131 , n5519 );
    not g28270 ( n8964 , n21293 );
    and g28271 ( n22130 , n19318 , n23670 );
    or g28272 ( n17747 , n17825 , n28107 );
    and g28273 ( n7259 , n6490 , n10958 );
    or g28274 ( n27567 , n18715 , n14402 );
    xnor g28275 ( n21339 , n26715 , n28948 );
    nor g28276 ( n23016 , n256 , n12285 );
    not g28277 ( n30988 , n27411 );
    xnor g28278 ( n26926 , n7315 , n29897 );
    or g28279 ( n20241 , n13834 , n27854 );
    not g28280 ( n5143 , n1575 );
    not g28281 ( n31659 , n547 );
    or g28282 ( n3230 , n30574 , n20832 );
    and g28283 ( n23295 , n31944 , n18163 );
    not g28284 ( n7307 , n10676 );
    and g28285 ( n24209 , n19446 , n20419 );
    not g28286 ( n6808 , n27452 );
    xnor g28287 ( n29424 , n30030 , n31528 );
    not g28288 ( n21003 , n16642 );
    not g28289 ( n25388 , n17772 );
    not g28290 ( n12990 , n3224 );
    nor g28291 ( n15622 , n534 , n28233 );
    or g28292 ( n16631 , n30398 , n18788 );
    xnor g28293 ( n30381 , n24713 , n2949 );
    nor g28294 ( n10124 , n26225 , n10557 );
    or g28295 ( n1938 , n12563 , n2111 );
    xnor g28296 ( n14932 , n31779 , n16227 );
    and g28297 ( n16272 , n18291 , n13716 );
    xor g28298 ( n12251 , n16697 , n3036 );
    not g28299 ( n4780 , n12159 );
    or g28300 ( n31747 , n9863 , n28037 );
    or g28301 ( n11170 , n12325 , n5690 );
    xnor g28302 ( n24789 , n21197 , n1954 );
    and g28303 ( n3479 , n12318 , n13796 );
    xnor g28304 ( n18352 , n25104 , n8345 );
    or g28305 ( n28841 , n4737 , n30978 );
    or g28306 ( n25222 , n3289 , n20981 );
    not g28307 ( n5229 , n28412 );
    and g28308 ( n23408 , n16700 , n12996 );
    or g28309 ( n9988 , n21186 , n30163 );
    not g28310 ( n10638 , n10879 );
    xnor g28311 ( n3985 , n5795 , n3290 );
    or g28312 ( n4823 , n8534 , n1743 );
    xnor g28313 ( n9918 , n25250 , n26379 );
    or g28314 ( n22542 , n21567 , n15177 );
    not g28315 ( n29017 , n12821 );
    nor g28316 ( n11328 , n26840 , n29011 );
    not g28317 ( n4047 , n24624 );
    xnor g28318 ( n30536 , n28760 , n23377 );
    or g28319 ( n10520 , n26257 , n22213 );
    not g28320 ( n7418 , n9816 );
    xnor g28321 ( n14471 , n23003 , n13454 );
    not g28322 ( n14496 , n10327 );
    nor g28323 ( n23684 , n27295 , n12118 );
    xnor g28324 ( n25559 , n4839 , n16425 );
    not g28325 ( n13831 , n8670 );
    and g28326 ( n15679 , n12670 , n7000 );
    or g28327 ( n7609 , n28517 , n28293 );
    and g28328 ( n10791 , n12436 , n23152 );
    or g28329 ( n30317 , n1115 , n30248 );
    xnor g28330 ( n16725 , n27034 , n29059 );
    not g28331 ( n30674 , n29187 );
    and g28332 ( n2715 , n11110 , n7638 );
    not g28333 ( n9289 , n19092 );
    xnor g28334 ( n18671 , n23877 , n1636 );
    xnor g28335 ( n24148 , n30732 , n21106 );
    or g28336 ( n21972 , n21140 , n13190 );
    xnor g28337 ( n26877 , n18948 , n8085 );
    not g28338 ( n23788 , n13157 );
    not g28339 ( n7316 , n5638 );
    or g28340 ( n26506 , n18319 , n14801 );
    and g28341 ( n16957 , n19732 , n9635 );
    not g28342 ( n12732 , n4133 );
    and g28343 ( n19726 , n22554 , n8498 );
    or g28344 ( n20702 , n14898 , n20229 );
    or g28345 ( n25634 , n6782 , n8039 );
    or g28346 ( n11525 , n3724 , n9463 );
    and g28347 ( n27049 , n16772 , n16149 );
    and g28348 ( n24560 , n14101 , n28048 );
    not g28349 ( n18453 , n31616 );
    not g28350 ( n16175 , n30105 );
    and g28351 ( n24145 , n13395 , n21469 );
    not g28352 ( n16891 , n19186 );
    or g28353 ( n6706 , n16595 , n26927 );
    xnor g28354 ( n11012 , n1110 , n24389 );
    xnor g28355 ( n6153 , n31673 , n29885 );
    not g28356 ( n393 , n25371 );
    not g28357 ( n11874 , n26491 );
    and g28358 ( n18186 , n18152 , n25967 );
    xnor g28359 ( n30390 , n20764 , n24131 );
    or g28360 ( n28093 , n22745 , n7376 );
    and g28361 ( n30886 , n10403 , n20221 );
    xnor g28362 ( n10565 , n3076 , n24429 );
    and g28363 ( n12516 , n20799 , n29090 );
    and g28364 ( n31538 , n3966 , n21920 );
    or g28365 ( n30168 , n16653 , n2513 );
    xor g28366 ( n2858 , n5744 , n20787 );
    or g28367 ( n12238 , n18706 , n25735 );
    and g28368 ( n15061 , n20500 , n25105 );
    or g28369 ( n7247 , n25378 , n11975 );
    or g28370 ( n23006 , n24902 , n15150 );
    xnor g28371 ( n30643 , n10332 , n11740 );
    xnor g28372 ( n18706 , n18934 , n18151 );
    not g28373 ( n6566 , n9670 );
    nor g28374 ( n22831 , n7143 , n26391 );
    not g28375 ( n11672 , n364 );
    or g28376 ( n28833 , n4187 , n15677 );
    xnor g28377 ( n27471 , n23461 , n3620 );
    or g28378 ( n30537 , n25334 , n19179 );
    xnor g28379 ( n8696 , n8454 , n28090 );
    and g28380 ( n22966 , n14935 , n10495 );
    not g28381 ( n13288 , n4450 );
    xnor g28382 ( n30502 , n4297 , n30536 );
    and g28383 ( n12622 , n15193 , n20648 );
    xnor g28384 ( n30445 , n13915 , n162 );
    and g28385 ( n2989 , n24360 , n28441 );
    xnor g28386 ( n27184 , n23847 , n6993 );
    and g28387 ( n4242 , n12541 , n23079 );
    not g28388 ( n10001 , n15035 );
    not g28389 ( n21316 , n27019 );
    or g28390 ( n13351 , n14187 , n8959 );
    not g28391 ( n24641 , n16639 );
    not g28392 ( n31120 , n18795 );
    xnor g28393 ( n13263 , n30457 , n23400 );
    or g28394 ( n18859 , n10136 , n13313 );
    or g28395 ( n12339 , n16901 , n14922 );
    xnor g28396 ( n28387 , n18667 , n8005 );
    and g28397 ( n16142 , n12359 , n3944 );
    or g28398 ( n9203 , n19032 , n13216 );
    nor g28399 ( n3635 , n25793 , n25613 );
    not g28400 ( n14492 , n233 );
    and g28401 ( n24411 , n26789 , n29394 );
    xnor g28402 ( n31139 , n12596 , n4632 );
    and g28403 ( n3499 , n10426 , n3706 );
    not g28404 ( n5193 , n22081 );
    xnor g28405 ( n22498 , n4125 , n2803 );
    xnor g28406 ( n3532 , n1840 , n27126 );
    or g28407 ( n17987 , n3806 , n30402 );
    xnor g28408 ( n21365 , n27666 , n7134 );
    and g28409 ( n26296 , n31294 , n13889 );
    and g28410 ( n29924 , n15498 , n9257 );
    xnor g28411 ( n19785 , n209 , n3440 );
    or g28412 ( n108 , n2610 , n29414 );
    xnor g28413 ( n2810 , n18394 , n16873 );
    or g28414 ( n28406 , n16787 , n7239 );
    xnor g28415 ( n4405 , n31169 , n3010 );
    and g28416 ( n31913 , n116 , n26389 );
    not g28417 ( n2830 , n16418 );
    or g28418 ( n7866 , n9460 , n12209 );
    nor g28419 ( n22269 , n22421 , n21015 );
    not g28420 ( n2326 , n5759 );
    or g28421 ( n3707 , n3364 , n29780 );
    not g28422 ( n4041 , n10029 );
    and g28423 ( n15973 , n9662 , n12590 );
    xnor g28424 ( n1823 , n28292 , n19892 );
    or g28425 ( n8442 , n19131 , n29160 );
    nor g28426 ( n1549 , n20600 , n28527 );
    or g28427 ( n11204 , n9948 , n8955 );
    and g28428 ( n27751 , n378 , n2602 );
    or g28429 ( n18050 , n10124 , n27098 );
    not g28430 ( n13913 , n1095 );
    not g28431 ( n23203 , n25028 );
    not g28432 ( n23207 , n26306 );
    and g28433 ( n20232 , n26267 , n12618 );
    and g28434 ( n28840 , n1271 , n4825 );
    or g28435 ( n538 , n11344 , n12344 );
    not g28436 ( n13502 , n29089 );
    not g28437 ( n13741 , n21133 );
    not g28438 ( n28247 , n22691 );
    xnor g28439 ( n26796 , n18975 , n7026 );
    or g28440 ( n22879 , n20416 , n9264 );
    not g28441 ( n23756 , n12401 );
    nor g28442 ( n13430 , n29568 , n9053 );
    or g28443 ( n29223 , n16379 , n4080 );
    not g28444 ( n20203 , n26828 );
    not g28445 ( n2928 , n21119 );
    nor g28446 ( n13096 , n21629 , n7022 );
    or g28447 ( n25901 , n30591 , n26309 );
    xnor g28448 ( n11920 , n11857 , n23151 );
    not g28449 ( n13978 , n24794 );
    nor g28450 ( n26344 , n15669 , n9792 );
    and g28451 ( n25354 , n4234 , n28128 );
    not g28452 ( n28555 , n13686 );
    not g28453 ( n12479 , n24807 );
    xnor g28454 ( n13451 , n28478 , n2062 );
    xnor g28455 ( n9259 , n23895 , n28713 );
    not g28456 ( n26252 , n15794 );
    and g28457 ( n27289 , n18456 , n31542 );
    not g28458 ( n21075 , n6273 );
    not g28459 ( n8526 , n21833 );
    or g28460 ( n21697 , n15396 , n15651 );
    or g28461 ( n9900 , n26327 , n18104 );
    xnor g28462 ( n5374 , n1874 , n30903 );
    not g28463 ( n25846 , n2728 );
    or g28464 ( n6821 , n8832 , n14218 );
    buf g28465 ( n29355 , n24490 );
    not g28466 ( n14573 , n27829 );
    not g28467 ( n21036 , n739 );
    xnor g28468 ( n22228 , n18761 , n4627 );
    not g28469 ( n20797 , n26410 );
    not g28470 ( n11974 , n23402 );
    not g28471 ( n5969 , n553 );
    not g28472 ( n4222 , n21822 );
    nor g28473 ( n20284 , n673 , n24940 );
    or g28474 ( n12789 , n29588 , n15070 );
    and g28475 ( n10986 , n4383 , n674 );
    or g28476 ( n25006 , n11112 , n5543 );
    xnor g28477 ( n6345 , n12566 , n891 );
    or g28478 ( n15872 , n4223 , n12801 );
    nor g28479 ( n25545 , n25616 , n8672 );
    xnor g28480 ( n28447 , n31260 , n21168 );
    or g28481 ( n21052 , n8888 , n29848 );
    xnor g28482 ( n2090 , n16119 , n13288 );
    not g28483 ( n22788 , n8732 );
    nor g28484 ( n11849 , n18380 , n13398 );
    or g28485 ( n30075 , n11308 , n21750 );
    or g28486 ( n18091 , n28299 , n31704 );
    xnor g28487 ( n17632 , n10698 , n20636 );
    xnor g28488 ( n23621 , n1097 , n7593 );
    xnor g28489 ( n9532 , n8728 , n20275 );
    or g28490 ( n10052 , n10737 , n22200 );
    nor g28491 ( n18009 , n21518 , n4941 );
    xnor g28492 ( n4057 , n16931 , n12352 );
    xnor g28493 ( n31233 , n3259 , n11736 );
    or g28494 ( n2125 , n751 , n19579 );
    buf g28495 ( n19003 , n20954 );
    not g28496 ( n29824 , n15485 );
    xnor g28497 ( n30984 , n10166 , n15369 );
    not g28498 ( n11705 , n7174 );
    and g28499 ( n26040 , n11199 , n27053 );
    or g28500 ( n10568 , n16267 , n27006 );
    not g28501 ( n25146 , n705 );
    or g28502 ( n23712 , n9243 , n26352 );
    not g28503 ( n29638 , n21784 );
    nor g28504 ( n25427 , n4662 , n30771 );
    or g28505 ( n25526 , n29472 , n8453 );
    not g28506 ( n30014 , n8584 );
    not g28507 ( n20051 , n25103 );
    xnor g28508 ( n22534 , n14823 , n16132 );
    or g28509 ( n8202 , n23313 , n10651 );
    not g28510 ( n12524 , n2629 );
    xnor g28511 ( n14695 , n18954 , n29375 );
    not g28512 ( n24418 , n18775 );
    and g28513 ( n15560 , n21594 , n24143 );
    or g28514 ( n1659 , n30950 , n15283 );
    xnor g28515 ( n3174 , n13642 , n21918 );
    nor g28516 ( n13423 , n1201 , n29921 );
    xnor g28517 ( n26466 , n11254 , n2210 );
    nor g28518 ( n23291 , n2319 , n7740 );
    nor g28519 ( n2833 , n30873 , n1767 );
    not g28520 ( n10397 , n24071 );
    or g28521 ( n21959 , n26356 , n29754 );
    or g28522 ( n1253 , n22868 , n2137 );
    and g28523 ( n9084 , n8148 , n14142 );
    or g28524 ( n8904 , n10964 , n10343 );
    and g28525 ( n8646 , n29446 , n16635 );
    or g28526 ( n22115 , n18376 , n7885 );
    xnor g28527 ( n11896 , n3776 , n29024 );
    or g28528 ( n21812 , n26338 , n23175 );
    or g28529 ( n13014 , n25083 , n5173 );
    or g28530 ( n29726 , n12451 , n251 );
    and g28531 ( n14170 , n26230 , n9013 );
    not g28532 ( n30983 , n29016 );
    and g28533 ( n24727 , n29951 , n29841 );
    or g28534 ( n18806 , n621 , n21068 );
    or g28535 ( n29219 , n30905 , n31112 );
    xnor g28536 ( n14835 , n7530 , n20235 );
    xnor g28537 ( n30624 , n7615 , n1515 );
    nor g28538 ( n28862 , n24132 , n30112 );
    not g28539 ( n8386 , n20871 );
    not g28540 ( n28920 , n22496 );
    and g28541 ( n5368 , n25935 , n3570 );
    or g28542 ( n24472 , n21382 , n3703 );
    and g28543 ( n2153 , n28351 , n21458 );
    not g28544 ( n13643 , n1027 );
    not g28545 ( n25330 , n16759 );
    nor g28546 ( n12108 , n16532 , n7149 );
    xnor g28547 ( n28472 , n445 , n5150 );
    or g28548 ( n23783 , n31086 , n12389 );
    xnor g28549 ( n11401 , n25240 , n4377 );
    nor g28550 ( n2148 , n15022 , n31942 );
    or g28551 ( n22132 , n4820 , n1814 );
    xnor g28552 ( n7903 , n3192 , n23203 );
    not g28553 ( n9645 , n236 );
    not g28554 ( n23876 , n23947 );
    xnor g28555 ( n17215 , n10617 , n29372 );
    xnor g28556 ( n15538 , n31953 , n13710 );
    xnor g28557 ( n18871 , n23612 , n27193 );
    or g28558 ( n20701 , n19412 , n3246 );
    and g28559 ( n30942 , n26152 , n14608 );
    or g28560 ( n23863 , n4963 , n3200 );
    not g28561 ( n18475 , n19965 );
    or g28562 ( n27942 , n29236 , n20595 );
    and g28563 ( n28971 , n4307 , n68 );
    xnor g28564 ( n18477 , n7414 , n14290 );
    xnor g28565 ( n26819 , n24086 , n9338 );
    not g28566 ( n17927 , n26061 );
    not g28567 ( n27379 , n31108 );
    not g28568 ( n31968 , n10785 );
    not g28569 ( n28571 , n7162 );
    and g28570 ( n5535 , n12752 , n24133 );
    nor g28571 ( n31179 , n24441 , n6320 );
    not g28572 ( n3682 , n16309 );
    xor g28573 ( n22958 , n8234 , n23306 );
    not g28574 ( n23158 , n9611 );
    and g28575 ( n20807 , n24930 , n15197 );
    not g28576 ( n21999 , n26002 );
    or g28577 ( n23793 , n12806 , n5108 );
    nor g28578 ( n1775 , n20388 , n721 );
    nor g28579 ( n2040 , n4648 , n25827 );
    or g28580 ( n27557 , n6446 , n18724 );
    xnor g28581 ( n10553 , n21095 , n11733 );
    xnor g28582 ( n21628 , n13824 , n20721 );
    and g28583 ( n25462 , n20264 , n28803 );
    nor g28584 ( n16026 , n31204 , n24769 );
    xnor g28585 ( n7965 , n6424 , n11169 );
    not g28586 ( n1527 , n8605 );
    or g28587 ( n14755 , n25106 , n10838 );
    nor g28588 ( n1269 , n13296 , n21951 );
    and g28589 ( n30016 , n30630 , n19141 );
    and g28590 ( n26760 , n249 , n30100 );
    nor g28591 ( n21056 , n2925 , n25805 );
    not g28592 ( n17548 , n30247 );
    and g28593 ( n11960 , n23881 , n17449 );
    and g28594 ( n19950 , n24390 , n7811 );
    not g28595 ( n30144 , n15020 );
    or g28596 ( n23981 , n3822 , n3688 );
    or g28597 ( n31899 , n17154 , n12326 );
    nor g28598 ( n17767 , n31595 , n11594 );
    or g28599 ( n9153 , n9948 , n21733 );
    and g28600 ( n15628 , n14190 , n10946 );
    and g28601 ( n8167 , n39 , n7238 );
    xnor g28602 ( n5392 , n5928 , n11689 );
    or g28603 ( n26779 , n10944 , n14190 );
    or g28604 ( n19884 , n12718 , n18520 );
    not g28605 ( n16912 , n28218 );
    and g28606 ( n27533 , n15721 , n11992 );
    xor g28607 ( n23740 , n26955 , n31973 );
    xnor g28608 ( n1637 , n3572 , n13137 );
    and g28609 ( n28513 , n32030 , n18634 );
    xnor g28610 ( n14854 , n28463 , n9377 );
    not g28611 ( n14317 , n5060 );
    or g28612 ( n7945 , n11462 , n16674 );
    xnor g28613 ( n3390 , n15615 , n5026 );
    not g28614 ( n21009 , n1702 );
    xnor g28615 ( n13849 , n11005 , n23789 );
    xnor g28616 ( n14779 , n2992 , n1713 );
    nor g28617 ( n19247 , n25889 , n12210 );
    not g28618 ( n19294 , n27969 );
    not g28619 ( n10241 , n26569 );
    not g28620 ( n131 , n17499 );
    or g28621 ( n27027 , n11789 , n6603 );
    xnor g28622 ( n5851 , n18667 , n19632 );
    xnor g28623 ( n13064 , n13272 , n4626 );
    xnor g28624 ( n22985 , n26156 , n10168 );
    and g28625 ( n19586 , n27892 , n3480 );
    not g28626 ( n6095 , n20341 );
    xnor g28627 ( n3999 , n23418 , n11692 );
    not g28628 ( n8077 , n31839 );
    not g28629 ( n7777 , n24066 );
    and g28630 ( n28554 , n31377 , n27338 );
    xnor g28631 ( n27452 , n30316 , n19388 );
    not g28632 ( n2232 , n25144 );
    or g28633 ( n6321 , n10756 , n13671 );
    and g28634 ( n27629 , n9922 , n5877 );
    xnor g28635 ( n14177 , n22045 , n6127 );
    and g28636 ( n29214 , n2699 , n19794 );
    not g28637 ( n17263 , n20274 );
    and g28638 ( n5502 , n14817 , n21943 );
    not g28639 ( n9754 , n29829 );
    not g28640 ( n7099 , n6726 );
    nor g28641 ( n1277 , n16019 , n3406 );
    xnor g28642 ( n27753 , n29615 , n18955 );
    or g28643 ( n18375 , n22320 , n18809 );
    xnor g28644 ( n20034 , n20781 , n5248 );
    and g28645 ( n9119 , n31364 , n12966 );
    not g28646 ( n2324 , n30411 );
    not g28647 ( n7248 , n28298 );
    xnor g28648 ( n17177 , n20738 , n7168 );
    and g28649 ( n15019 , n7599 , n8432 );
    or g28650 ( n22961 , n15847 , n11797 );
    or g28651 ( n21082 , n21210 , n15624 );
    not g28652 ( n5930 , n26284 );
    not g28653 ( n13242 , n27077 );
    or g28654 ( n15691 , n2237 , n15585 );
    and g28655 ( n13287 , n3277 , n1346 );
    not g28656 ( n28031 , n3255 );
    xnor g28657 ( n19873 , n16958 , n26867 );
    not g28658 ( n8813 , n2299 );
    xnor g28659 ( n17539 , n5696 , n29298 );
    xnor g28660 ( n16100 , n15588 , n30514 );
    not g28661 ( n29112 , n27955 );
    and g28662 ( n25110 , n3226 , n15875 );
    or g28663 ( n17277 , n8370 , n9134 );
    xnor g28664 ( n19843 , n27020 , n5045 );
    xnor g28665 ( n22548 , n22345 , n6888 );
    or g28666 ( n28455 , n30385 , n18348 );
    not g28667 ( n4813 , n11931 );
    or g28668 ( n32025 , n16873 , n27507 );
    not g28669 ( n18808 , n2610 );
    and g28670 ( n26546 , n10371 , n9813 );
    or g28671 ( n17532 , n9889 , n18031 );
    and g28672 ( n10750 , n27952 , n29375 );
    or g28673 ( n11369 , n28215 , n27515 );
    not g28674 ( n352 , n15748 );
    xnor g28675 ( n18230 , n6453 , n15219 );
    or g28676 ( n5943 , n2654 , n9129 );
    or g28677 ( n20162 , n16663 , n21578 );
    not g28678 ( n1855 , n11283 );
    xnor g28679 ( n17156 , n11364 , n17613 );
    xnor g28680 ( n12610 , n23688 , n12830 );
    not g28681 ( n5280 , n8804 );
    and g28682 ( n10698 , n7196 , n8047 );
    not g28683 ( n3959 , n12732 );
    xnor g28684 ( n7967 , n15513 , n10701 );
    and g28685 ( n934 , n23545 , n10778 );
    and g28686 ( n19840 , n18662 , n20150 );
    nor g28687 ( n2046 , n1616 , n30405 );
    or g28688 ( n30528 , n642 , n27975 );
    or g28689 ( n21001 , n9262 , n11679 );
    or g28690 ( n11639 , n5799 , n6050 );
    not g28691 ( n21679 , n4947 );
    xnor g28692 ( n31735 , n2553 , n23964 );
    nor g28693 ( n18262 , n11692 , n11116 );
    and g28694 ( n25143 , n23850 , n29427 );
    or g28695 ( n5495 , n3106 , n11244 );
    or g28696 ( n13163 , n16558 , n18496 );
    xnor g28697 ( n10825 , n14640 , n13423 );
    or g28698 ( n29287 , n1028 , n27063 );
    not g28699 ( n28250 , n2982 );
    xnor g28700 ( n4459 , n1627 , n8625 );
    xnor g28701 ( n25549 , n5873 , n18389 );
    or g28702 ( n12394 , n10509 , n31485 );
    or g28703 ( n15359 , n664 , n653 );
    xnor g28704 ( n2916 , n25046 , n6607 );
    not g28705 ( n3359 , n10550 );
    and g28706 ( n24606 , n28522 , n16647 );
    or g28707 ( n16669 , n19748 , n22891 );
    not g28708 ( n4981 , n16367 );
    not g28709 ( n8415 , n31000 );
    not g28710 ( n21212 , n25046 );
    and g28711 ( n16760 , n13739 , n23369 );
    xnor g28712 ( n13867 , n7201 , n9073 );
    or g28713 ( n25769 , n8474 , n9834 );
    or g28714 ( n22181 , n4860 , n26827 );
    or g28715 ( n15926 , n11835 , n5741 );
    not g28716 ( n22027 , n7220 );
    not g28717 ( n11352 , n25531 );
    not g28718 ( n26532 , n7025 );
    and g28719 ( n24869 , n10686 , n23169 );
    xnor g28720 ( n18684 , n20517 , n17019 );
    xnor g28721 ( n23615 , n3382 , n4524 );
    xor g28722 ( n31548 , n29414 , n698 );
    not g28723 ( n12817 , n24128 );
    xnor g28724 ( n14344 , n14735 , n2491 );
    or g28725 ( n31507 , n3214 , n5819 );
    or g28726 ( n18704 , n18586 , n27117 );
    not g28727 ( n14221 , n17460 );
    not g28728 ( n24920 , n21180 );
    xnor g28729 ( n31882 , n4655 , n8854 );
    or g28730 ( n20271 , n14345 , n14823 );
    or g28731 ( n18970 , n15788 , n6953 );
    not g28732 ( n26333 , n31881 );
    xnor g28733 ( n25441 , n31749 , n30213 );
    nor g28734 ( n21969 , n12892 , n12009 );
    not g28735 ( n18697 , n25569 );
    and g28736 ( n9668 , n10274 , n16846 );
    not g28737 ( n17511 , n9435 );
    nor g28738 ( n17508 , n20233 , n27538 );
    not g28739 ( n13985 , n20283 );
    or g28740 ( n27542 , n16113 , n12145 );
    and g28741 ( n25802 , n211 , n20245 );
    not g28742 ( n16281 , n17468 );
    or g28743 ( n5023 , n7647 , n20586 );
    not g28744 ( n364 , n27963 );
    nor g28745 ( n10732 , n27084 , n25374 );
    or g28746 ( n3899 , n27403 , n2698 );
    or g28747 ( n27712 , n21218 , n615 );
    nor g28748 ( n16901 , n7357 , n30597 );
    not g28749 ( n26200 , n12441 );
    or g28750 ( n26682 , n13536 , n3870 );
    xnor g28751 ( n21594 , n31530 , n21810 );
    xnor g28752 ( n17554 , n2786 , n25311 );
    and g28753 ( n8801 , n30551 , n5182 );
    or g28754 ( n4718 , n24477 , n1383 );
    not g28755 ( n8890 , n23980 );
    not g28756 ( n1767 , n6270 );
    not g28757 ( n4479 , n20552 );
    nor g28758 ( n9164 , n18735 , n21133 );
    nor g28759 ( n2951 , n22294 , n11016 );
    xnor g28760 ( n4680 , n23487 , n56 );
    xor g28761 ( n6480 , n26804 , n18086 );
    not g28762 ( n3531 , n3223 );
    xor g28763 ( n20764 , n12358 , n14852 );
    or g28764 ( n23021 , n14468 , n21742 );
    not g28765 ( n10109 , n23400 );
    or g28766 ( n5236 , n19820 , n17771 );
    xnor g28767 ( n16434 , n5081 , n17042 );
    and g28768 ( n9818 , n1894 , n31009 );
    xnor g28769 ( n10954 , n27998 , n3166 );
    not g28770 ( n18416 , n17126 );
    or g28771 ( n29903 , n15 , n3297 );
    not g28772 ( n25980 , n16998 );
    xnor g28773 ( n3728 , n19615 , n16406 );
    xnor g28774 ( n3169 , n7610 , n27880 );
    not g28775 ( n1333 , n12426 );
    and g28776 ( n18110 , n26322 , n1195 );
    xnor g28777 ( n12771 , n30407 , n31448 );
    xnor g28778 ( n11237 , n24325 , n30702 );
    and g28779 ( n26872 , n25294 , n14652 );
    xnor g28780 ( n15351 , n1076 , n31721 );
    not g28781 ( n21341 , n18164 );
    and g28782 ( n18291 , n2978 , n30660 );
    nor g28783 ( n9799 , n24429 , n11166 );
    and g28784 ( n13893 , n11939 , n6817 );
    not g28785 ( n21507 , n5905 );
    not g28786 ( n6140 , n20916 );
    or g28787 ( n14904 , n30456 , n28049 );
    or g28788 ( n24883 , n9588 , n26890 );
    or g28789 ( n25914 , n27080 , n15967 );
    not g28790 ( n12048 , n30758 );
    not g28791 ( n29294 , n434 );
    and g28792 ( n11263 , n17889 , n3211 );
    or g28793 ( n17228 , n13497 , n8842 );
    and g28794 ( n16267 , n20145 , n9882 );
    nor g28795 ( n15467 , n19194 , n7111 );
    xnor g28796 ( n26246 , n4771 , n27948 );
    and g28797 ( n12094 , n23425 , n25142 );
    and g28798 ( n29814 , n27840 , n11862 );
    nor g28799 ( n1754 , n21544 , n7535 );
    and g28800 ( n21602 , n5961 , n12362 );
    or g28801 ( n19530 , n7701 , n8124 );
    buf g28802 ( n29794 , n24795 );
    not g28803 ( n13330 , n21684 );
    and g28804 ( n31552 , n15814 , n14487 );
    not g28805 ( n5015 , n10413 );
    not g28806 ( n24834 , n2466 );
    nor g28807 ( n10924 , n793 , n23736 );
    xnor g28808 ( n28146 , n6509 , n31269 );
    not g28809 ( n10414 , n26502 );
    not g28810 ( n21933 , n20078 );
    or g28811 ( n2363 , n2371 , n934 );
    xnor g28812 ( n3775 , n3169 , n26365 );
    or g28813 ( n22873 , n14220 , n14692 );
    xnor g28814 ( n13105 , n4155 , n23591 );
    xnor g28815 ( n1280 , n16917 , n18402 );
    xnor g28816 ( n5942 , n534 , n20365 );
    not g28817 ( n17062 , n21697 );
    xnor g28818 ( n6056 , n13544 , n27768 );
    or g28819 ( n12420 , n22991 , n30507 );
    nor g28820 ( n21404 , n29444 , n24794 );
    or g28821 ( n29210 , n22151 , n27239 );
    xnor g28822 ( n14102 , n30488 , n25788 );
    not g28823 ( n17759 , n7677 );
    not g28824 ( n23622 , n24758 );
    not g28825 ( n17696 , n28180 );
    or g28826 ( n2380 , n14414 , n1576 );
    not g28827 ( n13370 , n7352 );
    xnor g28828 ( n30356 , n14723 , n31111 );
    not g28829 ( n2592 , n9744 );
    not g28830 ( n1137 , n26768 );
    and g28831 ( n20761 , n19711 , n18002 );
    or g28832 ( n10300 , n30328 , n7591 );
    nor g28833 ( n6324 , n10755 , n12280 );
    xnor g28834 ( n31362 , n26314 , n7688 );
    not g28835 ( n9759 , n19919 );
    and g28836 ( n30388 , n878 , n2940 );
    not g28837 ( n2872 , n16799 );
    or g28838 ( n7169 , n9133 , n16456 );
    xnor g28839 ( n24006 , n25929 , n12607 );
    and g28840 ( n31886 , n27665 , n82 );
    not g28841 ( n6816 , n2860 );
    or g28842 ( n13851 , n31787 , n8626 );
    and g28843 ( n9810 , n1594 , n11329 );
    and g28844 ( n12822 , n12369 , n27794 );
    and g28845 ( n27644 , n15571 , n30058 );
    or g28846 ( n23351 , n6626 , n22405 );
    not g28847 ( n3780 , n1461 );
    or g28848 ( n18888 , n31610 , n11786 );
    and g28849 ( n27522 , n17885 , n26368 );
    nor g28850 ( n20409 , n25069 , n12597 );
    nor g28851 ( n2470 , n23770 , n10430 );
    xnor g28852 ( n20160 , n31414 , n17851 );
    or g28853 ( n8136 , n4654 , n27415 );
    or g28854 ( n30548 , n13254 , n22251 );
    or g28855 ( n17944 , n637 , n5554 );
    xnor g28856 ( n7030 , n7978 , n12143 );
    or g28857 ( n6795 , n13189 , n26503 );
    and g28858 ( n9015 , n1058 , n24644 );
    or g28859 ( n20083 , n4048 , n30858 );
    xnor g28860 ( n9873 , n22359 , n30811 );
    or g28861 ( n15729 , n29733 , n13674 );
    not g28862 ( n2943 , n4735 );
    not g28863 ( n2744 , n775 );
    xnor g28864 ( n15511 , n7750 , n11891 );
    and g28865 ( n5465 , n22786 , n11637 );
    and g28866 ( n6214 , n26311 , n2480 );
    not g28867 ( n16385 , n27041 );
    not g28868 ( n9892 , n15311 );
    or g28869 ( n5676 , n6352 , n14346 );
    or g28870 ( n8982 , n22550 , n18562 );
    not g28871 ( n31976 , n28468 );
    not g28872 ( n12664 , n17305 );
    and g28873 ( n774 , n7483 , n8786 );
    or g28874 ( n3801 , n22209 , n12622 );
    nor g28875 ( n14588 , n24070 , n20603 );
    and g28876 ( n9814 , n5589 , n17577 );
    not g28877 ( n12280 , n30426 );
    and g28878 ( n26740 , n4823 , n26570 );
    xnor g28879 ( n14802 , n8829 , n15293 );
    xnor g28880 ( n26062 , n2483 , n18955 );
    not g28881 ( n8188 , n12597 );
    or g28882 ( n24904 , n757 , n4946 );
    and g28883 ( n16761 , n18978 , n19656 );
    or g28884 ( n30987 , n14763 , n1334 );
    or g28885 ( n2612 , n8371 , n20752 );
    and g28886 ( n28538 , n22833 , n21538 );
    xnor g28887 ( n30042 , n29754 , n7801 );
    not g28888 ( n4210 , n12118 );
    xnor g28889 ( n7862 , n20405 , n11402 );
    not g28890 ( n22634 , n17184 );
    or g28891 ( n14028 , n9423 , n9887 );
    and g28892 ( n14367 , n2580 , n10215 );
    nor g28893 ( n1372 , n28376 , n31954 );
    or g28894 ( n28176 , n23136 , n10328 );
    not g28895 ( n25525 , n26552 );
    or g28896 ( n19390 , n4607 , n8327 );
    xnor g28897 ( n30318 , n18323 , n15944 );
    xnor g28898 ( n28963 , n7794 , n24598 );
    xnor g28899 ( n15027 , n11164 , n24717 );
    not g28900 ( n22635 , n25880 );
    or g28901 ( n24348 , n3924 , n14885 );
    not g28902 ( n15170 , n12486 );
    and g28903 ( n17078 , n9232 , n10894 );
    and g28904 ( n2636 , n20111 , n368 );
    not g28905 ( n11239 , n13259 );
    and g28906 ( n31791 , n28707 , n12815 );
    and g28907 ( n17399 , n25751 , n28461 );
    xnor g28908 ( n29883 , n26506 , n31830 );
    or g28909 ( n15594 , n5788 , n29857 );
    or g28910 ( n19451 , n31407 , n30860 );
    xnor g28911 ( n18690 , n272 , n608 );
    xnor g28912 ( n13472 , n7108 , n19035 );
    and g28913 ( n27740 , n3155 , n28782 );
    and g28914 ( n13337 , n10719 , n17114 );
    or g28915 ( n12985 , n16840 , n26736 );
    and g28916 ( n6622 , n27604 , n27124 );
    xor g28917 ( n10627 , n23321 , n29897 );
    xnor g28918 ( n16104 , n12881 , n16610 );
    or g28919 ( n30196 , n12952 , n21789 );
    xnor g28920 ( n16415 , n26859 , n10893 );
    and g28921 ( n3941 , n24339 , n23318 );
    or g28922 ( n28728 , n3173 , n31033 );
    nor g28923 ( n31920 , n7359 , n952 );
    xnor g28924 ( n23655 , n27623 , n2204 );
    xnor g28925 ( n22395 , n12614 , n9474 );
    or g28926 ( n31642 , n4818 , n21388 );
    xnor g28927 ( n19847 , n20113 , n15993 );
    xnor g28928 ( n7161 , n5104 , n17715 );
    or g28929 ( n10618 , n12721 , n9018 );
    nor g28930 ( n23245 , n22176 , n10489 );
    not g28931 ( n11138 , n22935 );
    and g28932 ( n22439 , n24845 , n30241 );
    not g28933 ( n2811 , n26974 );
    or g28934 ( n28284 , n8089 , n8154 );
    xnor g28935 ( n19979 , n3260 , n26375 );
    and g28936 ( n15206 , n15200 , n11696 );
    or g28937 ( n22074 , n22139 , n20451 );
    not g28938 ( n22331 , n9469 );
    nor g28939 ( n5856 , n31481 , n17429 );
    xnor g28940 ( n30846 , n11320 , n16389 );
    xnor g28941 ( n402 , n13475 , n9239 );
    not g28942 ( n26258 , n9601 );
    not g28943 ( n7531 , n10323 );
    xnor g28944 ( n16427 , n7259 , n28303 );
    xnor g28945 ( n3653 , n30619 , n27904 );
    not g28946 ( n26182 , n9478 );
    xnor g28947 ( n26080 , n16075 , n30201 );
    and g28948 ( n2957 , n1956 , n6436 );
    and g28949 ( n18430 , n1456 , n23186 );
    nor g28950 ( n19330 , n23117 , n27609 );
    or g28951 ( n628 , n30468 , n20587 );
    or g28952 ( n1364 , n11853 , n19351 );
    and g28953 ( n185 , n31568 , n15118 );
    or g28954 ( n14673 , n15301 , n14268 );
    nor g28955 ( n29786 , n5559 , n27535 );
    not g28956 ( n29673 , n18189 );
    and g28957 ( n31400 , n29894 , n9050 );
    or g28958 ( n26614 , n6306 , n17561 );
    or g28959 ( n8569 , n8142 , n15916 );
    or g28960 ( n26010 , n29850 , n19682 );
    xnor g28961 ( n4863 , n15738 , n14214 );
    or g28962 ( n5002 , n2571 , n131 );
    xnor g28963 ( n18153 , n9721 , n4799 );
    not g28964 ( n22626 , n2340 );
    and g28965 ( n11291 , n9047 , n20826 );
    or g28966 ( n28995 , n6125 , n17118 );
    and g28967 ( n31900 , n13721 , n31602 );
    not g28968 ( n8250 , n3333 );
    or g28969 ( n24058 , n29249 , n1302 );
    not g28970 ( n4397 , n20961 );
    and g28971 ( n20674 , n25106 , n20293 );
    not g28972 ( n7219 , n5523 );
    and g28973 ( n23452 , n539 , n7906 );
    not g28974 ( n29172 , n4556 );
    not g28975 ( n24990 , n4531 );
    or g28976 ( n24375 , n27235 , n13436 );
    xnor g28977 ( n3781 , n7180 , n5783 );
    xnor g28978 ( n14024 , n18843 , n10207 );
    nor g28979 ( n24285 , n15366 , n7734 );
    not g28980 ( n3117 , n10056 );
    or g28981 ( n11020 , n13020 , n2103 );
    not g28982 ( n15052 , n22111 );
    or g28983 ( n7139 , n209 , n3595 );
    or g28984 ( n23228 , n1616 , n10563 );
    not g28985 ( n30882 , n29673 );
    xnor g28986 ( n31493 , n30306 , n32009 );
    or g28987 ( n3384 , n29112 , n25472 );
    not g28988 ( n31176 , n5674 );
    not g28989 ( n3362 , n26541 );
    or g28990 ( n18123 , n4538 , n11787 );
    not g28991 ( n20 , n8822 );
    or g28992 ( n11292 , n29401 , n17076 );
    xor g28993 ( n16287 , n30491 , n256 );
    not g28994 ( n11918 , n21803 );
    or g28995 ( n9212 , n16821 , n16360 );
    xnor g28996 ( n19883 , n22303 , n23443 );
    and g28997 ( n2250 , n3073 , n5862 );
    or g28998 ( n26457 , n28150 , n14546 );
    xnor g28999 ( n14615 , n19378 , n6422 );
    or g29000 ( n7972 , n26953 , n11476 );
    not g29001 ( n6257 , n555 );
    xnor g29002 ( n9774 , n17216 , n8133 );
    not g29003 ( n22844 , n4644 );
    nor g29004 ( n14117 , n20038 , n5879 );
    or g29005 ( n5269 , n6223 , n1010 );
    xnor g29006 ( n27959 , n664 , n17255 );
    or g29007 ( n11329 , n10196 , n25157 );
    not g29008 ( n24573 , n9751 );
    not g29009 ( n16356 , n4434 );
    or g29010 ( n10297 , n24525 , n23957 );
    and g29011 ( n27862 , n7790 , n31064 );
    not g29012 ( n20471 , n6944 );
    or g29013 ( n24237 , n31623 , n456 );
    and g29014 ( n17352 , n12106 , n11986 );
    or g29015 ( n12270 , n8530 , n19213 );
    and g29016 ( n2057 , n25363 , n23917 );
    not g29017 ( n18509 , n11981 );
    nor g29018 ( n20532 , n21034 , n840 );
    or g29019 ( n25840 , n1545 , n4696 );
    or g29020 ( n8350 , n28011 , n5509 );
    nor g29021 ( n28023 , n24304 , n5599 );
    or g29022 ( n31550 , n24504 , n10791 );
    xnor g29023 ( n30797 , n13567 , n15050 );
    not g29024 ( n24149 , n1304 );
    or g29025 ( n28473 , n23268 , n12631 );
    or g29026 ( n6793 , n8573 , n15186 );
    and g29027 ( n30979 , n21095 , n18213 );
    xnor g29028 ( n26854 , n19874 , n14503 );
    or g29029 ( n16781 , n16654 , n9754 );
    xnor g29030 ( n4819 , n28861 , n12895 );
    xnor g29031 ( n23357 , n19066 , n24712 );
    xnor g29032 ( n11128 , n16803 , n23342 );
    and g29033 ( n20217 , n17535 , n12818 );
    xnor g29034 ( n23539 , n15105 , n9321 );
    not g29035 ( n8963 , n10451 );
    not g29036 ( n18572 , n1202 );
    xor g29037 ( n19107 , n9821 , n17970 );
    xnor g29038 ( n17416 , n13214 , n21355 );
    not g29039 ( n5730 , n20341 );
    nor g29040 ( n28174 , n2520 , n5101 );
    xnor g29041 ( n3567 , n14692 , n14272 );
    xnor g29042 ( n18151 , n3830 , n26786 );
    or g29043 ( n5648 , n9464 , n22424 );
    not g29044 ( n8881 , n13326 );
    not g29045 ( n3919 , n2535 );
    xnor g29046 ( n8567 , n25704 , n4393 );
    not g29047 ( n25000 , n5675 );
    not g29048 ( n29616 , n8613 );
    not g29049 ( n12097 , n12634 );
    or g29050 ( n26570 , n21161 , n7672 );
    or g29051 ( n14803 , n9335 , n18494 );
    or g29052 ( n9577 , n31142 , n8607 );
    not g29053 ( n30122 , n16637 );
    xnor g29054 ( n23395 , n7559 , n4335 );
    or g29055 ( n5681 , n31572 , n27066 );
    and g29056 ( n50 , n4178 , n11449 );
    xnor g29057 ( n854 , n10425 , n6981 );
    not g29058 ( n14021 , n29307 );
    or g29059 ( n27265 , n497 , n15704 );
    not g29060 ( n19513 , n18691 );
    not g29061 ( n5123 , n10222 );
    nor g29062 ( n13039 , n14558 , n22053 );
    or g29063 ( n3754 , n6122 , n14734 );
    xnor g29064 ( n4503 , n3966 , n2605 );
    or g29065 ( n1627 , n6148 , n24641 );
    not g29066 ( n17753 , n3124 );
    and g29067 ( n11000 , n6644 , n17961 );
    nor g29068 ( n25215 , n25579 , n17729 );
    and g29069 ( n13508 , n25796 , n22434 );
    or g29070 ( n10086 , n30381 , n2524 );
    xnor g29071 ( n24651 , n31462 , n5715 );
    not g29072 ( n27523 , n20015 );
    not g29073 ( n13343 , n24578 );
    not g29074 ( n14506 , n29202 );
    not g29075 ( n721 , n14324 );
    or g29076 ( n1090 , n22819 , n31126 );
    xnor g29077 ( n24242 , n19404 , n29355 );
    nor g29078 ( n15877 , n25431 , n8694 );
    xnor g29079 ( n17651 , n21554 , n31344 );
    nor g29080 ( n5316 , n3259 , n11736 );
    or g29081 ( n21501 , n4001 , n24751 );
    not g29082 ( n12815 , n20052 );
    xnor g29083 ( n20986 , n17252 , n26297 );
    and g29084 ( n16380 , n12606 , n10003 );
    not g29085 ( n18804 , n5684 );
    not g29086 ( n29930 , n22059 );
    xnor g29087 ( n27562 , n26519 , n6543 );
    not g29088 ( n16848 , n22296 );
    not g29089 ( n17533 , n31474 );
    xnor g29090 ( n6469 , n10814 , n9486 );
    xnor g29091 ( n30606 , n20167 , n28058 );
    nor g29092 ( n20157 , n1057 , n10802 );
    xnor g29093 ( n6204 , n12935 , n26581 );
    not g29094 ( n28213 , n8478 );
    nor g29095 ( n17639 , n3649 , n2853 );
    or g29096 ( n10217 , n7287 , n13091 );
    nor g29097 ( n8315 , n25365 , n12009 );
    not g29098 ( n6060 , n25793 );
    not g29099 ( n3058 , n13723 );
    nor g29100 ( n11371 , n12288 , n26717 );
    xnor g29101 ( n7198 , n15303 , n6309 );
    or g29102 ( n25005 , n21785 , n9938 );
    xnor g29103 ( n6915 , n6393 , n6372 );
    nor g29104 ( n12968 , n3814 , n17389 );
    and g29105 ( n11726 , n9602 , n25712 );
    or g29106 ( n5595 , n31708 , n18926 );
    xnor g29107 ( n17768 , n4706 , n17830 );
    xnor g29108 ( n27601 , n6333 , n23319 );
    xnor g29109 ( n15840 , n14233 , n2798 );
    xnor g29110 ( n11550 , n13677 , n18002 );
    not g29111 ( n15830 , n27416 );
    and g29112 ( n5375 , n9683 , n18518 );
    or g29113 ( n24073 , n17019 , n11394 );
    not g29114 ( n4007 , n708 );
    not g29115 ( n24323 , n8710 );
    xnor g29116 ( n15465 , n13852 , n22942 );
    not g29117 ( n1971 , n15917 );
    or g29118 ( n26649 , n5905 , n3689 );
    or g29119 ( n16351 , n29435 , n29785 );
    nor g29120 ( n11951 , n25430 , n22781 );
    or g29121 ( n2893 , n28274 , n7673 );
    or g29122 ( n4842 , n7184 , n7943 );
    nor g29123 ( n18041 , n19960 , n9931 );
    not g29124 ( n20428 , n17108 );
    and g29125 ( n4672 , n12203 , n28774 );
    not g29126 ( n272 , n4451 );
    or g29127 ( n16405 , n20208 , n15810 );
    and g29128 ( n15554 , n21576 , n9230 );
    nor g29129 ( n19263 , n15135 , n31681 );
    not g29130 ( n567 , n29553 );
    xnor g29131 ( n28231 , n30191 , n17677 );
    nor g29132 ( n28605 , n1196 , n4284 );
    xnor g29133 ( n9258 , n2035 , n13239 );
    or g29134 ( n10337 , n23795 , n31825 );
    not g29135 ( n25646 , n24525 );
    and g29136 ( n19024 , n794 , n20535 );
    xnor g29137 ( n16382 , n13322 , n24028 );
    xnor g29138 ( n26960 , n17392 , n16545 );
    not g29139 ( n335 , n3002 );
    not g29140 ( n22637 , n8592 );
    and g29141 ( n15685 , n755 , n30868 );
    not g29142 ( n13885 , n24049 );
    or g29143 ( n15984 , n20122 , n21627 );
    or g29144 ( n28964 , n24392 , n27995 );
    or g29145 ( n1758 , n13314 , n23265 );
    xnor g29146 ( n19913 , n16761 , n12623 );
    or g29147 ( n5427 , n10937 , n15721 );
    or g29148 ( n30197 , n10895 , n6597 );
    and g29149 ( n2572 , n16016 , n16992 );
    xnor g29150 ( n13389 , n5129 , n7532 );
    or g29151 ( n17266 , n28010 , n1240 );
    xnor g29152 ( n3778 , n25357 , n7640 );
    not g29153 ( n19288 , n19920 );
    not g29154 ( n19311 , n16174 );
    or g29155 ( n11687 , n21057 , n6840 );
    xnor g29156 ( n6291 , n18667 , n30405 );
    xnor g29157 ( n8797 , n2515 , n16558 );
    and g29158 ( n29872 , n30451 , n31040 );
    and g29159 ( n15871 , n7296 , n4704 );
    or g29160 ( n20813 , n22015 , n21620 );
    and g29161 ( n5590 , n8105 , n25185 );
    or g29162 ( n3871 , n29215 , n22507 );
    not g29163 ( n10871 , n13790 );
    xnor g29164 ( n31057 , n10107 , n10455 );
    xnor g29165 ( n28786 , n27340 , n20563 );
    xnor g29166 ( n28311 , n12888 , n25495 );
    xnor g29167 ( n30367 , n20442 , n11711 );
    or g29168 ( n3868 , n8645 , n7806 );
    not g29169 ( n32016 , n21321 );
    xnor g29170 ( n26410 , n6285 , n20448 );
    and g29171 ( n20893 , n15747 , n564 );
    nor g29172 ( n8431 , n26894 , n23966 );
    not g29173 ( n7546 , n133 );
    and g29174 ( n22083 , n1968 , n12337 );
    or g29175 ( n4565 , n7528 , n5808 );
    nor g29176 ( n26870 , n6916 , n24116 );
    xnor g29177 ( n14141 , n25760 , n3268 );
    xnor g29178 ( n28281 , n4537 , n24194 );
    nor g29179 ( n22706 , n775 , n29798 );
    nor g29180 ( n7567 , n8263 , n27941 );
    not g29181 ( n2105 , n9745 );
    and g29182 ( n7181 , n10644 , n11084 );
    xnor g29183 ( n21138 , n7981 , n5561 );
    or g29184 ( n16265 , n31147 , n7530 );
    xnor g29185 ( n28622 , n2985 , n16872 );
    not g29186 ( n1036 , n30343 );
    and g29187 ( n18014 , n8921 , n13241 );
    not g29188 ( n23463 , n24783 );
    not g29189 ( n22551 , n30754 );
    or g29190 ( n9470 , n14925 , n9578 );
    not g29191 ( n4828 , n4490 );
    or g29192 ( n10329 , n22717 , n22836 );
    xnor g29193 ( n31789 , n18476 , n11233 );
    not g29194 ( n32028 , n479 );
    not g29195 ( n20474 , n21961 );
    not g29196 ( n15598 , n1039 );
    xnor g29197 ( n13301 , n11122 , n1165 );
    xnor g29198 ( n17015 , n3307 , n20799 );
    not g29199 ( n30867 , n29932 );
    or g29200 ( n5606 , n8705 , n18915 );
    xnor g29201 ( n2631 , n20834 , n26724 );
    xnor g29202 ( n21754 , n27947 , n31066 );
    xnor g29203 ( n12972 , n18507 , n28634 );
    or g29204 ( n4431 , n3996 , n20865 );
    xnor g29205 ( n74 , n23096 , n13756 );
    not g29206 ( n19054 , n6940 );
    xnor g29207 ( n9978 , n1346 , n28180 );
    or g29208 ( n27465 , n1635 , n2408 );
    not g29209 ( n2640 , n21954 );
    and g29210 ( n4761 , n1121 , n11243 );
    and g29211 ( n3502 , n9986 , n30386 );
    and g29212 ( n14364 , n15235 , n13936 );
    not g29213 ( n19801 , n21748 );
    xnor g29214 ( n12158 , n8724 , n28772 );
    and g29215 ( n10285 , n18123 , n24461 );
    nor g29216 ( n10469 , n26929 , n3745 );
    xnor g29217 ( n28543 , n13107 , n20904 );
    and g29218 ( n17157 , n29272 , n1887 );
    xnor g29219 ( n23979 , n9480 , n18475 );
    or g29220 ( n13386 , n30251 , n22876 );
    and g29221 ( n9679 , n25926 , n10981 );
    not g29222 ( n4556 , n21208 );
    not g29223 ( n4311 , n2146 );
    not g29224 ( n28365 , n23772 );
    xnor g29225 ( n22632 , n9101 , n24210 );
    or g29226 ( n5466 , n14310 , n23447 );
    not g29227 ( n28545 , n29739 );
    xnor g29228 ( n2528 , n4390 , n27030 );
    and g29229 ( n27287 , n17005 , n24371 );
    and g29230 ( n28789 , n22422 , n17089 );
    not g29231 ( n6974 , n17298 );
    and g29232 ( n7149 , n9784 , n1114 );
    not g29233 ( n10624 , n18918 );
    not g29234 ( n2677 , n4898 );
    xnor g29235 ( n9254 , n18391 , n27233 );
    nor g29236 ( n4362 , n11218 , n21384 );
    and g29237 ( n1286 , n12403 , n3481 );
    xnor g29238 ( n28899 , n23320 , n24289 );
    not g29239 ( n18180 , n8710 );
    xnor g29240 ( n5 , n19012 , n9159 );
    xor g29241 ( n481 , n19328 , n21185 );
    and g29242 ( n16572 , n25135 , n21019 );
    xnor g29243 ( n6137 , n4340 , n14984 );
    nor g29244 ( n21271 , n28616 , n21248 );
    not g29245 ( n20861 , n30346 );
    not g29246 ( n10973 , n3313 );
    not g29247 ( n31961 , n3545 );
    buf g29248 ( n16583 , n30124 );
    and g29249 ( n21857 , n3300 , n22727 );
    or g29250 ( n12239 , n7051 , n28237 );
    xnor g29251 ( n36 , n25982 , n4554 );
    nor g29252 ( n30558 , n23956 , n26331 );
    or g29253 ( n28457 , n22095 , n3002 );
    xor g29254 ( n15857 , n5176 , n17650 );
    and g29255 ( n14733 , n7079 , n10998 );
    xnor g29256 ( n5635 , n10490 , n12024 );
    and g29257 ( n18056 , n27543 , n10195 );
    xor g29258 ( n11837 , n26066 , n9679 );
    buf g29259 ( n26029 , n105 );
    nor g29260 ( n17179 , n11526 , n2603 );
    not g29261 ( n18595 , n14503 );
    xor g29262 ( n5255 , n19729 , n8711 );
    not g29263 ( n29948 , n26525 );
    not g29264 ( n23912 , n22470 );
    or g29265 ( n10500 , n19310 , n28119 );
    not g29266 ( n24976 , n23605 );
    or g29267 ( n25067 , n17381 , n19961 );
    xnor g29268 ( n18139 , n25921 , n21530 );
    or g29269 ( n17500 , n21271 , n15089 );
    not g29270 ( n9527 , n1404 );
    and g29271 ( n12029 , n17897 , n8823 );
    not g29272 ( n22384 , n18829 );
    xnor g29273 ( n16494 , n10435 , n8392 );
    and g29274 ( n20364 , n16506 , n26759 );
    not g29275 ( n24647 , n26255 );
    or g29276 ( n8653 , n29020 , n13311 );
    or g29277 ( n19296 , n3550 , n3961 );
    and g29278 ( n8877 , n23085 , n13133 );
    and g29279 ( n10020 , n4008 , n27803 );
    not g29280 ( n7778 , n2866 );
    or g29281 ( n7914 , n3144 , n5794 );
    nor g29282 ( n25008 , n27595 , n19788 );
    not g29283 ( n21648 , n21034 );
    and g29284 ( n909 , n29817 , n22408 );
    not g29285 ( n17132 , n10301 );
    xor g29286 ( n29019 , n2048 , n3534 );
    or g29287 ( n8096 , n3025 , n17757 );
    not g29288 ( n23903 , n23365 );
    and g29289 ( n21627 , n3476 , n7782 );
    not g29290 ( n22928 , n5378 );
    not g29291 ( n2948 , n28920 );
    not g29292 ( n26005 , n12649 );
    xnor g29293 ( n30801 , n14299 , n15976 );
    or g29294 ( n29113 , n6423 , n27115 );
    not g29295 ( n27521 , n5753 );
    and g29296 ( n9184 , n18422 , n20461 );
    not g29297 ( n27498 , n24595 );
    and g29298 ( n2710 , n12365 , n25312 );
    not g29299 ( n2742 , n28797 );
    not g29300 ( n25708 , n24137 );
    and g29301 ( n27811 , n11604 , n16995 );
    nor g29302 ( n31567 , n20890 , n7723 );
    not g29303 ( n23839 , n26387 );
    or g29304 ( n9196 , n13312 , n7412 );
    not g29305 ( n20629 , n18419 );
    xor g29306 ( n11215 , n12058 , n24557 );
    nor g29307 ( n14676 , n12566 , n25653 );
    not g29308 ( n11290 , n24569 );
    and g29309 ( n10390 , n3456 , n15594 );
    nor g29310 ( n9583 , n25242 , n24122 );
    nor g29311 ( n8645 , n18165 , n27154 );
    or g29312 ( n29800 , n29639 , n8930 );
    xor g29313 ( n17386 , n2196 , n27170 );
    xnor g29314 ( n14426 , n31563 , n19817 );
    not g29315 ( n7909 , n3569 );
    or g29316 ( n26099 , n17013 , n19749 );
    not g29317 ( n2033 , n13003 );
    and g29318 ( n30779 , n29616 , n5029 );
    not g29319 ( n17440 , n27500 );
    not g29320 ( n5091 , n17226 );
    not g29321 ( n27743 , n12433 );
    or g29322 ( n19436 , n12542 , n7879 );
    or g29323 ( n13755 , n4081 , n14321 );
    and g29324 ( n29928 , n17410 , n29048 );
    xnor g29325 ( n21813 , n3222 , n12687 );
    xnor g29326 ( n30432 , n18160 , n19987 );
    not g29327 ( n13625 , n4604 );
    or g29328 ( n4870 , n26769 , n29970 );
    xnor g29329 ( n3105 , n12906 , n30723 );
    xnor g29330 ( n1091 , n26175 , n19881 );
    or g29331 ( n9448 , n20578 , n4755 );
    and g29332 ( n25153 , n22785 , n11061 );
    or g29333 ( n7628 , n6296 , n55 );
    not g29334 ( n10559 , n18706 );
    not g29335 ( n11044 , n20052 );
    xnor g29336 ( n26381 , n30409 , n24879 );
    xnor g29337 ( n6365 , n26015 , n18112 );
    not g29338 ( n18651 , n31417 );
    and g29339 ( n6652 , n16677 , n18489 );
    or g29340 ( n25671 , n5089 , n31709 );
    or g29341 ( n25785 , n24397 , n6392 );
    xnor g29342 ( n23902 , n18402 , n28376 );
    and g29343 ( n1576 , n7119 , n11898 );
    not g29344 ( n18561 , n27002 );
    xnor g29345 ( n8676 , n5834 , n4278 );
    xnor g29346 ( n15783 , n22916 , n2520 );
    xnor g29347 ( n15271 , n14759 , n15336 );
    xnor g29348 ( n22902 , n3721 , n23317 );
    xnor g29349 ( n9822 , n15 , n23218 );
    or g29350 ( n5366 , n4723 , n24365 );
    nor g29351 ( n24699 , n24414 , n3443 );
    not g29352 ( n29898 , n4188 );
    xnor g29353 ( n30719 , n7593 , n9338 );
    not g29354 ( n11287 , n1543 );
    and g29355 ( n15437 , n19875 , n13080 );
    or g29356 ( n26079 , n28956 , n20863 );
    and g29357 ( n14575 , n7737 , n12792 );
    and g29358 ( n31995 , n31156 , n25218 );
    or g29359 ( n14619 , n28369 , n9868 );
    or g29360 ( n8086 , n26082 , n6060 );
    and g29361 ( n183 , n5207 , n25039 );
    not g29362 ( n28112 , n5319 );
    not g29363 ( n24094 , n23871 );
    not g29364 ( n10181 , n27461 );
    not g29365 ( n19458 , n28396 );
    nor g29366 ( n4352 , n15152 , n12867 );
    not g29367 ( n22842 , n32021 );
    and g29368 ( n2782 , n7484 , n6996 );
    xnor g29369 ( n2156 , n27275 , n8210 );
    or g29370 ( n28895 , n11836 , n26264 );
    not g29371 ( n2918 , n9680 );
    xnor g29372 ( n4771 , n10387 , n660 );
    not g29373 ( n20357 , n13067 );
    and g29374 ( n16697 , n20306 , n13172 );
    or g29375 ( n31657 , n31718 , n4995 );
    and g29376 ( n4974 , n14786 , n22807 );
    not g29377 ( n16428 , n74 );
    or g29378 ( n17490 , n2230 , n29852 );
    xnor g29379 ( n5893 , n15506 , n21730 );
    xnor g29380 ( n17468 , n18811 , n29859 );
    or g29381 ( n10033 , n8229 , n14130 );
    xnor g29382 ( n3936 , n10765 , n16229 );
    not g29383 ( n24975 , n7539 );
    not g29384 ( n31992 , n19312 );
    not g29385 ( n1886 , n11319 );
    or g29386 ( n16877 , n7359 , n24653 );
    nor g29387 ( n20142 , n8133 , n17216 );
    xnor g29388 ( n11743 , n12837 , n15396 );
    and g29389 ( n17070 , n2125 , n31922 );
    xnor g29390 ( n5580 , n26646 , n4505 );
    xnor g29391 ( n23135 , n23879 , n397 );
    xnor g29392 ( n20730 , n16860 , n7258 );
    xnor g29393 ( n2291 , n12800 , n17385 );
    not g29394 ( n24029 , n7762 );
    nor g29395 ( n14187 , n15762 , n8347 );
    and g29396 ( n15459 , n4337 , n10089 );
    or g29397 ( n24847 , n10102 , n29071 );
    xnor g29398 ( n2433 , n10788 , n21549 );
    not g29399 ( n31957 , n729 );
    xnor g29400 ( n26007 , n19039 , n29195 );
    xnor g29401 ( n5073 , n16841 , n6976 );
    xnor g29402 ( n12726 , n13426 , n28622 );
    and g29403 ( n2639 , n21951 , n27956 );
    xnor g29404 ( n22197 , n11669 , n13843 );
    xnor g29405 ( n28796 , n14539 , n22345 );
    not g29406 ( n27786 , n26130 );
    or g29407 ( n11351 , n8963 , n23279 );
    nor g29408 ( n7711 , n18412 , n13268 );
    xnor g29409 ( n30789 , n11100 , n16540 );
    and g29410 ( n3316 , n10189 , n20061 );
    xnor g29411 ( n30165 , n23008 , n418 );
    xnor g29412 ( n9670 , n9905 , n24971 );
    and g29413 ( n14897 , n18708 , n25129 );
    not g29414 ( n28896 , n8670 );
    not g29415 ( n8972 , n27334 );
    and g29416 ( n31142 , n29922 , n10549 );
    not g29417 ( n14292 , n25999 );
    nor g29418 ( n10509 , n16112 , n5276 );
    or g29419 ( n20661 , n22379 , n7109 );
    xnor g29420 ( n31428 , n8381 , n23047 );
    and g29421 ( n23658 , n24950 , n31238 );
    nor g29422 ( n14633 , n11658 , n16609 );
    or g29423 ( n5815 , n10414 , n3913 );
    or g29424 ( n26703 , n11360 , n24365 );
    xnor g29425 ( n22385 , n19983 , n26867 );
    not g29426 ( n21800 , n9999 );
    or g29427 ( n7058 , n21804 , n6077 );
    or g29428 ( n28181 , n25032 , n9222 );
    xnor g29429 ( n7588 , n17113 , n25490 );
    and g29430 ( n31687 , n24393 , n31597 );
    xnor g29431 ( n5112 , n11130 , n15678 );
    not g29432 ( n19378 , n7204 );
    xnor g29433 ( n20562 , n15361 , n21310 );
    or g29434 ( n22365 , n29575 , n22001 );
    or g29435 ( n30737 , n20715 , n7071 );
    not g29436 ( n11712 , n29527 );
    xnor g29437 ( n367 , n24118 , n2798 );
    not g29438 ( n1027 , n21677 );
    or g29439 ( n4548 , n20630 , n947 );
    or g29440 ( n22426 , n10954 , n30992 );
    xnor g29441 ( n29733 , n696 , n3009 );
    and g29442 ( n22544 , n30574 , n20691 );
    not g29443 ( n9040 , n3299 );
    and g29444 ( n28005 , n1897 , n27590 );
    or g29445 ( n2590 , n9965 , n11557 );
    not g29446 ( n5260 , n14962 );
    or g29447 ( n10121 , n23205 , n9190 );
    nor g29448 ( n1282 , n5388 , n25206 );
    xnor g29449 ( n2059 , n17511 , n26668 );
    xnor g29450 ( n29076 , n13977 , n18033 );
    not g29451 ( n12036 , n8558 );
    not g29452 ( n22377 , n18577 );
    xnor g29453 ( n7879 , n14913 , n12591 );
    or g29454 ( n23545 , n25828 , n2130 );
    or g29455 ( n2795 , n29347 , n243 );
    xnor g29456 ( n25577 , n15269 , n445 );
    xnor g29457 ( n19289 , n13751 , n15382 );
    or g29458 ( n7000 , n30887 , n25063 );
    or g29459 ( n14832 , n14204 , n19395 );
    not g29460 ( n18929 , n13287 );
    nor g29461 ( n25939 , n16806 , n20427 );
    not g29462 ( n30103 , n18331 );
    and g29463 ( n12646 , n4021 , n20206 );
    and g29464 ( n573 , n28236 , n790 );
    and g29465 ( n16564 , n5035 , n27576 );
    or g29466 ( n5926 , n26911 , n8219 );
    and g29467 ( n29716 , n4126 , n12528 );
    or g29468 ( n14075 , n31980 , n6678 );
    xnor g29469 ( n12922 , n5600 , n24530 );
    or g29470 ( n30734 , n23402 , n6305 );
    not g29471 ( n24852 , n31868 );
    not g29472 ( n3631 , n22866 );
    or g29473 ( n19580 , n17227 , n21771 );
    or g29474 ( n13459 , n747 , n4632 );
    or g29475 ( n23830 , n25881 , n28740 );
    not g29476 ( n17775 , n9783 );
    not g29477 ( n7458 , n5485 );
    not g29478 ( n19711 , n434 );
    or g29479 ( n11832 , n16640 , n12176 );
    or g29480 ( n2387 , n8941 , n21729 );
    xnor g29481 ( n20998 , n4831 , n5439 );
    and g29482 ( n19854 , n9170 , n1739 );
    and g29483 ( n11808 , n28439 , n27263 );
    and g29484 ( n15264 , n6073 , n12447 );
    xnor g29485 ( n22960 , n30078 , n18702 );
    and g29486 ( n13458 , n29099 , n10372 );
    or g29487 ( n25752 , n23291 , n6479 );
    or g29488 ( n19568 , n17735 , n29753 );
    and g29489 ( n11551 , n29300 , n28972 );
    or g29490 ( n7773 , n12853 , n134 );
    xnor g29491 ( n14197 , n135 , n17146 );
    or g29492 ( n16850 , n24345 , n20743 );
    not g29493 ( n8763 , n11886 );
    not g29494 ( n11348 , n1151 );
    not g29495 ( n17479 , n21950 );
    buf g29496 ( n15272 , n10699 );
    xnor g29497 ( n30703 , n30001 , n3478 );
    not g29498 ( n16524 , n4877 );
    and g29499 ( n10441 , n15217 , n8438 );
    or g29500 ( n19608 , n1764 , n30864 );
    not g29501 ( n3142 , n15156 );
    or g29502 ( n25905 , n14182 , n24815 );
    not g29503 ( n26559 , n17111 );
    not g29504 ( n23853 , n7213 );
    or g29505 ( n20694 , n7060 , n16212 );
    or g29506 ( n10318 , n17598 , n17789 );
    not g29507 ( n4526 , n12781 );
    and g29508 ( n7974 , n18296 , n16364 );
    xnor g29509 ( n19280 , n9780 , n525 );
    not g29510 ( n17903 , n9569 );
    not g29511 ( n28369 , n12179 );
    xnor g29512 ( n12830 , n6016 , n18177 );
    or g29513 ( n8744 , n21372 , n5479 );
    not g29514 ( n12079 , n16312 );
    or g29515 ( n26448 , n11047 , n19256 );
    xnor g29516 ( n6558 , n13987 , n10350 );
    and g29517 ( n4502 , n17608 , n12386 );
    and g29518 ( n28424 , n14664 , n8759 );
    and g29519 ( n22877 , n10092 , n21185 );
    xnor g29520 ( n4933 , n16700 , n27365 );
    not g29521 ( n19747 , n17257 );
    xnor g29522 ( n24478 , n23625 , n11411 );
    or g29523 ( n7008 , n27284 , n21325 );
    xnor g29524 ( n5371 , n14951 , n24536 );
    not g29525 ( n10735 , n20704 );
    and g29526 ( n18044 , n7846 , n9916 );
    not g29527 ( n7021 , n11037 );
    or g29528 ( n8604 , n22244 , n6322 );
    or g29529 ( n10258 , n25524 , n3524 );
    or g29530 ( n14048 , n24956 , n28886 );
    xnor g29531 ( n23899 , n30229 , n15299 );
    xnor g29532 ( n31380 , n21919 , n20739 );
    not g29533 ( n16687 , n31391 );
    or g29534 ( n15841 , n10158 , n4274 );
    or g29535 ( n7066 , n31669 , n14245 );
    or g29536 ( n26201 , n341 , n25855 );
    nor g29537 ( n28915 , n3396 , n6401 );
    not g29538 ( n5136 , n6873 );
    or g29539 ( n13353 , n20079 , n11673 );
    xnor g29540 ( n22367 , n20605 , n19334 );
    or g29541 ( n94 , n4983 , n5609 );
    not g29542 ( n19363 , n21909 );
    not g29543 ( n5037 , n9317 );
    xnor g29544 ( n2053 , n4461 , n2655 );
    not g29545 ( n18843 , n1856 );
    not g29546 ( n29557 , n15771 );
    or g29547 ( n5678 , n19493 , n12308 );
    not g29548 ( n17331 , n6651 );
    xnor g29549 ( n19959 , n482 , n843 );
    xnor g29550 ( n22855 , n4470 , n20495 );
    or g29551 ( n19286 , n4345 , n28933 );
    nor g29552 ( n1468 , n6682 , n31749 );
    xnor g29553 ( n6813 , n1470 , n16093 );
    nor g29554 ( n7034 , n11120 , n6474 );
    not g29555 ( n8909 , n7675 );
    not g29556 ( n22904 , n26487 );
    xnor g29557 ( n16024 , n24611 , n8702 );
    or g29558 ( n1362 , n12511 , n4435 );
    xnor g29559 ( n15322 , n24548 , n3683 );
    xnor g29560 ( n14613 , n8205 , n17170 );
    not g29561 ( n1719 , n10420 );
    xnor g29562 ( n22455 , n6917 , n24118 );
    or g29563 ( n14115 , n24090 , n17393 );
    not g29564 ( n27831 , n7751 );
    or g29565 ( n20426 , n22208 , n15655 );
    xnor g29566 ( n7044 , n354 , n22719 );
    and g29567 ( n1173 , n12296 , n7699 );
    and g29568 ( n30859 , n26672 , n7837 );
    nor g29569 ( n5116 , n27316 , n28390 );
    and g29570 ( n2919 , n2882 , n13275 );
    nor g29571 ( n21807 , n16131 , n31007 );
    and g29572 ( n1743 , n2692 , n16497 );
    nor g29573 ( n6177 , n12379 , n6068 );
    not g29574 ( n10073 , n4404 );
    xnor g29575 ( n16545 , n17915 , n5066 );
    not g29576 ( n18583 , n28044 );
    xnor g29577 ( n16252 , n23661 , n14666 );
    xnor g29578 ( n13619 , n194 , n12746 );
    not g29579 ( n4240 , n16711 );
    or g29580 ( n2310 , n6111 , n27538 );
    xor g29581 ( n18296 , n16639 , n3828 );
    xnor g29582 ( n5261 , n31274 , n599 );
    buf g29583 ( n16660 , n17672 );
    xnor g29584 ( n22302 , n2444 , n21186 );
    not g29585 ( n3404 , n2669 );
    not g29586 ( n29262 , n16587 );
    or g29587 ( n16486 , n173 , n11872 );
    xnor g29588 ( n13936 , n18556 , n18477 );
    not g29589 ( n26202 , n27883 );
    nor g29590 ( n21657 , n27021 , n28502 );
    and g29591 ( n3099 , n16988 , n1123 );
    buf g29592 ( n2453 , n6487 );
    or g29593 ( n27306 , n28072 , n8769 );
    and g29594 ( n26725 , n27294 , n17679 );
    not g29595 ( n10468 , n25953 );
    not g29596 ( n27253 , n8152 );
    or g29597 ( n19063 , n9297 , n7652 );
    or g29598 ( n20912 , n17101 , n8830 );
    xnor g29599 ( n30004 , n14971 , n5851 );
    not g29600 ( n16864 , n25204 );
    and g29601 ( n7134 , n12698 , n15139 );
    and g29602 ( n29500 , n13402 , n8014 );
    or g29603 ( n2575 , n2609 , n10986 );
    xnor g29604 ( n15126 , n27233 , n15436 );
    not g29605 ( n13292 , n18645 );
    not g29606 ( n17983 , n5873 );
    or g29607 ( n24109 , n14697 , n3053 );
    or g29608 ( n12792 , n11265 , n17963 );
    nor g29609 ( n8275 , n3782 , n27354 );
    or g29610 ( n19230 , n3785 , n8467 );
    or g29611 ( n26701 , n29669 , n30563 );
    not g29612 ( n13124 , n26505 );
    xnor g29613 ( n30678 , n12368 , n3754 );
    xnor g29614 ( n11997 , n3205 , n28663 );
    or g29615 ( n29202 , n28676 , n1734 );
    not g29616 ( n4201 , n16002 );
    not g29617 ( n11579 , n7180 );
    xnor g29618 ( n7801 , n23379 , n800 );
    not g29619 ( n25971 , n27253 );
    xnor g29620 ( n23255 , n23337 , n17899 );
    not g29621 ( n17220 , n24525 );
    or g29622 ( n19509 , n27832 , n30208 );
    not g29623 ( n24221 , n4973 );
    and g29624 ( n7835 , n19296 , n2523 );
    not g29625 ( n22372 , n24926 );
    and g29626 ( n2080 , n23913 , n8810 );
    not g29627 ( n17036 , n30201 );
    not g29628 ( n27876 , n6865 );
    or g29629 ( n21917 , n23097 , n12573 );
    and g29630 ( n8707 , n9888 , n22643 );
    not g29631 ( n20663 , n8333 );
    xnor g29632 ( n20603 , n28120 , n10882 );
    not g29633 ( n14147 , n18429 );
    or g29634 ( n30406 , n10451 , n25514 );
    not g29635 ( n4561 , n16267 );
    not g29636 ( n20253 , n10185 );
    nor g29637 ( n21230 , n14962 , n14333 );
    not g29638 ( n29297 , n21882 );
    and g29639 ( n31729 , n21514 , n8901 );
    xnor g29640 ( n25891 , n10188 , n17150 );
    or g29641 ( n20163 , n16994 , n27146 );
    or g29642 ( n5154 , n29702 , n24049 );
    not g29643 ( n25389 , n2137 );
    not g29644 ( n17200 , n26624 );
    xnor g29645 ( n27405 , n29581 , n16783 );
    xnor g29646 ( n13819 , n12315 , n18830 );
    nor g29647 ( n17158 , n632 , n12364 );
    or g29648 ( n13030 , n31367 , n15885 );
    xnor g29649 ( n2330 , n11836 , n30458 );
    not g29650 ( n7892 , n8774 );
    or g29651 ( n1969 , n12552 , n24033 );
    or g29652 ( n8730 , n1498 , n16854 );
    not g29653 ( n27147 , n10071 );
    xnor g29654 ( n14469 , n22930 , n29550 );
    or g29655 ( n5904 , n2384 , n7467 );
    not g29656 ( n17757 , n15674 );
    nor g29657 ( n7861 , n30831 , n2539 );
    or g29658 ( n6891 , n21000 , n21877 );
    and g29659 ( n24035 , n18360 , n22665 );
    not g29660 ( n19600 , n26743 );
    not g29661 ( n10869 , n18874 );
    or g29662 ( n14727 , n11643 , n25646 );
    or g29663 ( n6906 , n5312 , n5405 );
    nor g29664 ( n16757 , n25422 , n7283 );
    not g29665 ( n6003 , n959 );
    not g29666 ( n9615 , n2086 );
    xnor g29667 ( n16216 , n6882 , n16075 );
    xnor g29668 ( n22929 , n27907 , n18685 );
    not g29669 ( n28950 , n9803 );
    or g29670 ( n13805 , n11296 , n5909 );
    nor g29671 ( n29639 , n13318 , n8173 );
    not g29672 ( n1934 , n129 );
    not g29673 ( n19464 , n24464 );
    xnor g29674 ( n11651 , n23733 , n3121 );
    or g29675 ( n7949 , n15014 , n26157 );
    xnor g29676 ( n6304 , n25334 , n19231 );
    and g29677 ( n11675 , n27481 , n11468 );
    and g29678 ( n23301 , n23113 , n11769 );
    and g29679 ( n2482 , n10593 , n23882 );
    or g29680 ( n19635 , n27255 , n11977 );
    nor g29681 ( n3836 , n3307 , n28736 );
    and g29682 ( n20479 , n31779 , n3989 );
    and g29683 ( n23683 , n30623 , n1450 );
    not g29684 ( n21829 , n26191 );
    not g29685 ( n14894 , n6974 );
    not g29686 ( n2519 , n4003 );
    and g29687 ( n19353 , n26044 , n6007 );
    xnor g29688 ( n27407 , n5695 , n22550 );
    or g29689 ( n22627 , n14702 , n1168 );
    xnor g29690 ( n5243 , n31444 , n6291 );
    or g29691 ( n25118 , n9330 , n6907 );
    or g29692 ( n20580 , n8546 , n4575 );
    xnor g29693 ( n8715 , n27916 , n24584 );
    not g29694 ( n29912 , n24289 );
    or g29695 ( n17608 , n15862 , n28579 );
    and g29696 ( n225 , n11012 , n735 );
    xnor g29697 ( n525 , n15833 , n31595 );
    buf g29698 ( n17090 , n125 );
    xnor g29699 ( n5215 , n6673 , n18387 );
    not g29700 ( n31420 , n20365 );
    not g29701 ( n908 , n9776 );
    xnor g29702 ( n12715 , n21261 , n22867 );
    not g29703 ( n26256 , n23978 );
    xnor g29704 ( n18985 , n864 , n20467 );
    and g29705 ( n1768 , n6350 , n20726 );
    and g29706 ( n19414 , n27593 , n8204 );
    or g29707 ( n25672 , n10711 , n3761 );
    or g29708 ( n21118 , n12588 , n23180 );
    not g29709 ( n17226 , n3702 );
    xnor g29710 ( n21994 , n5663 , n8611 );
    xnor g29711 ( n21215 , n7319 , n30823 );
    nor g29712 ( n25806 , n17797 , n30029 );
    not g29713 ( n437 , n27352 );
    not g29714 ( n22659 , n30525 );
    xnor g29715 ( n5766 , n12030 , n9655 );
    and g29716 ( n13622 , n29985 , n28553 );
    nor g29717 ( n12647 , n6626 , n3968 );
    or g29718 ( n12913 , n28873 , n26407 );
    and g29719 ( n16211 , n29518 , n27350 );
    or g29720 ( n9348 , n20210 , n8503 );
    xnor g29721 ( n18570 , n7587 , n1057 );
    xnor g29722 ( n6180 , n7517 , n18460 );
    not g29723 ( n12634 , n5867 );
    not g29724 ( n17971 , n18296 );
    xnor g29725 ( n1325 , n20705 , n15364 );
    or g29726 ( n22658 , n21111 , n4868 );
    not g29727 ( n5768 , n28611 );
    xnor g29728 ( n24783 , n8793 , n11531 );
    xnor g29729 ( n23444 , n20363 , n20183 );
    not g29730 ( n8122 , n20345 );
    and g29731 ( n5309 , n15420 , n30017 );
    not g29732 ( n4865 , n27459 );
    or g29733 ( n11213 , n20761 , n28371 );
    or g29734 ( n14749 , n20497 , n104 );
    or g29735 ( n5167 , n21004 , n29755 );
    xnor g29736 ( n799 , n9726 , n16709 );
    not g29737 ( n11965 , n4086 );
    and g29738 ( n30595 , n9794 , n21995 );
    or g29739 ( n10704 , n30481 , n25200 );
    or g29740 ( n21053 , n16756 , n5677 );
    not g29741 ( n17389 , n29971 );
    not g29742 ( n16006 , n16559 );
    and g29743 ( n32033 , n19449 , n18925 );
    not g29744 ( n11387 , n6885 );
    or g29745 ( n31209 , n1055 , n8669 );
    xnor g29746 ( n8064 , n16715 , n19435 );
    xnor g29747 ( n24575 , n28729 , n24612 );
    not g29748 ( n2555 , n8713 );
    xnor g29749 ( n467 , n13140 , n28815 );
    not g29750 ( n28756 , n20917 );
    xnor g29751 ( n11655 , n30039 , n5742 );
    xnor g29752 ( n5448 , n19790 , n17499 );
    xnor g29753 ( n5661 , n11751 , n13230 );
    and g29754 ( n31075 , n337 , n10579 );
    or g29755 ( n4689 , n15588 , n30514 );
    xnor g29756 ( n13876 , n1199 , n7431 );
    nor g29757 ( n201 , n16633 , n24440 );
    or g29758 ( n10415 , n2981 , n10068 );
    or g29759 ( n14293 , n7593 , n6243 );
    and g29760 ( n26954 , n29191 , n11463 );
    not g29761 ( n23292 , n5588 );
    or g29762 ( n2752 , n10751 , n16832 );
    not g29763 ( n5752 , n16132 );
    and g29764 ( n7823 , n1822 , n24927 );
    not g29765 ( n1769 , n24858 );
    or g29766 ( n20867 , n26060 , n31362 );
    or g29767 ( n15990 , n31497 , n23844 );
    not g29768 ( n15638 , n7184 );
    not g29769 ( n16978 , n13976 );
    nor g29770 ( n28986 , n27574 , n513 );
    or g29771 ( n7097 , n20534 , n5790 );
    nor g29772 ( n3339 , n6681 , n30339 );
    not g29773 ( n18960 , n31689 );
    not g29774 ( n9910 , n11712 );
    or g29775 ( n18185 , n3162 , n28005 );
    or g29776 ( n17560 , n31923 , n8780 );
    not g29777 ( n22919 , n20726 );
    xnor g29778 ( n26858 , n21268 , n4684 );
    not g29779 ( n16177 , n10477 );
    and g29780 ( n1941 , n14805 , n14489 );
    or g29781 ( n14877 , n19370 , n11417 );
    not g29782 ( n212 , n21212 );
    or g29783 ( n2426 , n22671 , n19491 );
    or g29784 ( n2393 , n16944 , n617 );
    or g29785 ( n165 , n9799 , n22018 );
    nor g29786 ( n14096 , n18394 , n30334 );
    xnor g29787 ( n2340 , n20652 , n462 );
    not g29788 ( n22390 , n31566 );
    not g29789 ( n25013 , n29840 );
    not g29790 ( n30090 , n2512 );
    and g29791 ( n12995 , n5364 , n9082 );
    nor g29792 ( n14859 , n10847 , n3422 );
    xnor g29793 ( n27978 , n23735 , n2963 );
    or g29794 ( n26671 , n30343 , n22399 );
    or g29795 ( n24692 , n14661 , n10362 );
    or g29796 ( n4364 , n26188 , n15770 );
    xnor g29797 ( n13560 , n7494 , n15964 );
    not g29798 ( n21410 , n21901 );
    or g29799 ( n17450 , n10556 , n13481 );
    xnor g29800 ( n18267 , n2948 , n2564 );
    or g29801 ( n24746 , n11421 , n11901 );
    and g29802 ( n10432 , n23257 , n21134 );
    not g29803 ( n8844 , n16746 );
    or g29804 ( n15474 , n21482 , n1183 );
    nor g29805 ( n19098 , n21597 , n19000 );
    not g29806 ( n14410 , n10049 );
    and g29807 ( n16408 , n23848 , n28634 );
    not g29808 ( n27276 , n26179 );
    and g29809 ( n2042 , n2795 , n23589 );
    not g29810 ( n19862 , n15408 );
    xnor g29811 ( n28788 , n31142 , n1096 );
    not g29812 ( n4092 , n9104 );
    xnor g29813 ( n9752 , n25889 , n12210 );
    xnor g29814 ( n25502 , n5860 , n22134 );
    and g29815 ( n24183 , n23093 , n21770 );
    and g29816 ( n21641 , n5429 , n28900 );
    not g29817 ( n3799 , n3992 );
    xnor g29818 ( n21767 , n18222 , n18684 );
    not g29819 ( n12900 , n14940 );
    or g29820 ( n15193 , n29500 , n5702 );
    or g29821 ( n29742 , n28577 , n13626 );
    not g29822 ( n30199 , n26584 );
    xnor g29823 ( n25190 , n28402 , n27002 );
    and g29824 ( n17603 , n2497 , n7863 );
    nor g29825 ( n4200 , n4748 , n21037 );
    or g29826 ( n14639 , n3863 , n14185 );
    not g29827 ( n1590 , n27534 );
    not g29828 ( n14566 , n3106 );
    not g29829 ( n2430 , n14915 );
    or g29830 ( n22097 , n7951 , n27345 );
    nor g29831 ( n7164 , n18547 , n17565 );
    not g29832 ( n19357 , n3021 );
    xnor g29833 ( n21673 , n28737 , n12625 );
    xnor g29834 ( n16053 , n18285 , n20518 );
    nor g29835 ( n14176 , n7046 , n12443 );
    and g29836 ( n22625 , n7560 , n9336 );
    nor g29837 ( n13447 , n20121 , n18366 );
    not g29838 ( n29952 , n15311 );
    and g29839 ( n6457 , n31834 , n25617 );
    or g29840 ( n4380 , n11717 , n22027 );
    not g29841 ( n14255 , n23359 );
    and g29842 ( n8196 , n13342 , n22156 );
    or g29843 ( n26053 , n21818 , n25547 );
    and g29844 ( n10679 , n8405 , n6764 );
    xnor g29845 ( n4641 , n18286 , n31918 );
    xnor g29846 ( n28870 , n21555 , n769 );
    or g29847 ( n12321 , n4138 , n8131 );
    or g29848 ( n7114 , n16525 , n23037 );
    not g29849 ( n14772 , n26212 );
    or g29850 ( n9813 , n31573 , n18832 );
    not g29851 ( n5323 , n14298 );
    xnor g29852 ( n6039 , n1034 , n796 );
    and g29853 ( n6834 , n8036 , n15893 );
    not g29854 ( n13726 , n9625 );
    or g29855 ( n29504 , n8476 , n19040 );
    xnor g29856 ( n28131 , n14444 , n9060 );
    nor g29857 ( n13773 , n1720 , n16304 );
    xnor g29858 ( n5511 , n21715 , n24187 );
    xnor g29859 ( n10040 , n14007 , n22656 );
    nor g29860 ( n7570 , n12618 , n13431 );
    or g29861 ( n26310 , n29355 , n18936 );
    xnor g29862 ( n10839 , n15308 , n4533 );
    not g29863 ( n18617 , n9241 );
    xnor g29864 ( n3733 , n29032 , n20630 );
    not g29865 ( n13232 , n17233 );
    xnor g29866 ( n15453 , n15718 , n3166 );
    or g29867 ( n25340 , n12753 , n21287 );
    or g29868 ( n21285 , n28012 , n12702 );
    and g29869 ( n16236 , n16244 , n4069 );
    and g29870 ( n28544 , n25916 , n6561 );
    not g29871 ( n30491 , n26261 );
    xnor g29872 ( n31915 , n27931 , n19762 );
    not g29873 ( n6637 , n5642 );
    or g29874 ( n26431 , n6636 , n60 );
    not g29875 ( n23122 , n20475 );
    and g29876 ( n11968 , n10702 , n24731 );
    xnor g29877 ( n10447 , n8573 , n11868 );
    not g29878 ( n8531 , n20913 );
    or g29879 ( n11604 , n15324 , n23048 );
    not g29880 ( n31379 , n12425 );
    or g29881 ( n30675 , n23898 , n20029 );
    and g29882 ( n7375 , n23367 , n7269 );
    not g29883 ( n1119 , n23340 );
    nor g29884 ( n14204 , n21135 , n29363 );
    not g29885 ( n16014 , n23588 );
    and g29886 ( n20010 , n30644 , n247 );
    not g29887 ( n9865 , n1507 );
    not g29888 ( n11385 , n7768 );
    and g29889 ( n8044 , n9442 , n11877 );
    xnor g29890 ( n12511 , n2131 , n26809 );
    nor g29891 ( n9777 , n22858 , n18820 );
    xnor g29892 ( n7943 , n9870 , n15028 );
    nor g29893 ( n15082 , n15363 , n20041 );
    or g29894 ( n29404 , n30562 , n19887 );
    xnor g29895 ( n17194 , n15117 , n18878 );
    and g29896 ( n22435 , n15660 , n12548 );
    or g29897 ( n3379 , n23865 , n8812 );
    xnor g29898 ( n3774 , n10433 , n30201 );
    and g29899 ( n8179 , n15327 , n16622 );
    and g29900 ( n8039 , n10465 , n10972 );
    not g29901 ( n17599 , n26346 );
    xnor g29902 ( n3951 , n22098 , n13372 );
    and g29903 ( n27068 , n14700 , n30139 );
    xnor g29904 ( n1018 , n15704 , n22766 );
    xnor g29905 ( n8928 , n102 , n30028 );
    xnor g29906 ( n8223 , n20799 , n2939 );
    xnor g29907 ( n13841 , n13301 , n11740 );
    or g29908 ( n10915 , n31710 , n18300 );
    xnor g29909 ( n11379 , n8919 , n3036 );
    or g29910 ( n18635 , n22602 , n5249 );
    not g29911 ( n3223 , n14135 );
    and g29912 ( n3125 , n10625 , n28641 );
    or g29913 ( n15388 , n16498 , n29281 );
    xor g29914 ( n303 , n17038 , n24794 );
    not g29915 ( n21589 , n23596 );
    or g29916 ( n7483 , n6389 , n29096 );
    or g29917 ( n30372 , n12240 , n17777 );
    not g29918 ( n29645 , n6168 );
    xnor g29919 ( n27830 , n3735 , n23910 );
    and g29920 ( n2266 , n24562 , n22476 );
    not g29921 ( n30636 , n7770 );
    not g29922 ( n13852 , n2791 );
    xnor g29923 ( n26878 , n9011 , n14112 );
    not g29924 ( n29397 , n15999 );
    not g29925 ( n1304 , n7154 );
    not g29926 ( n13491 , n15849 );
    not g29927 ( n28194 , n29615 );
    xnor g29928 ( n5298 , n1177 , n20038 );
    or g29929 ( n19539 , n31788 , n4691 );
    nor g29930 ( n2274 , n14227 , n19092 );
    and g29931 ( n22461 , n30542 , n22297 );
    or g29932 ( n15907 , n17003 , n8946 );
    and g29933 ( n31262 , n2958 , n25862 );
    and g29934 ( n17728 , n20758 , n25141 );
    and g29935 ( n2650 , n4462 , n6567 );
    not g29936 ( n6708 , n2836 );
    not g29937 ( n20982 , n28787 );
    xnor g29938 ( n10943 , n691 , n25966 );
    not g29939 ( n21087 , n29016 );
    and g29940 ( n9035 , n11817 , n6045 );
    not g29941 ( n5284 , n21647 );
    not g29942 ( n443 , n31481 );
    xnor g29943 ( n18758 , n19943 , n4130 );
    nor g29944 ( n8045 , n28734 , n4246 );
    nor g29945 ( n18632 , n28233 , n7378 );
    not g29946 ( n26067 , n2354 );
    xnor g29947 ( n9561 , n17140 , n3489 );
    not g29948 ( n966 , n27210 );
    xnor g29949 ( n19011 , n4216 , n20535 );
    or g29950 ( n11326 , n12786 , n20924 );
    and g29951 ( n30183 , n7739 , n15389 );
    and g29952 ( n30912 , n30462 , n7049 );
    nor g29953 ( n31596 , n17125 , n3401 );
    or g29954 ( n13943 , n8472 , n19661 );
    or g29955 ( n6774 , n18922 , n18260 );
    not g29956 ( n28590 , n26403 );
    or g29957 ( n2819 , n30825 , n14776 );
    or g29958 ( n11126 , n18696 , n27872 );
    xnor g29959 ( n8485 , n23977 , n919 );
    not g29960 ( n1107 , n14489 );
    xnor g29961 ( n2847 , n14358 , n6779 );
    or g29962 ( n20693 , n22967 , n2406 );
    xnor g29963 ( n27594 , n29685 , n17633 );
    not g29964 ( n29798 , n21585 );
    or g29965 ( n8923 , n10093 , n13093 );
    or g29966 ( n19499 , n16162 , n13794 );
    xnor g29967 ( n17828 , n197 , n5188 );
    not g29968 ( n11423 , n15847 );
    not g29969 ( n23095 , n17952 );
    xnor g29970 ( n11101 , n31541 , n31590 );
    not g29971 ( n10259 , n18955 );
    not g29972 ( n28559 , n23769 );
    xnor g29973 ( n21529 , n12597 , n9239 );
    and g29974 ( n26318 , n3362 , n6603 );
    or g29975 ( n25244 , n10287 , n5596 );
    xnor g29976 ( n8939 , n5450 , n20874 );
    and g29977 ( n26635 , n30007 , n31329 );
    not g29978 ( n24662 , n24239 );
    not g29979 ( n5114 , n3251 );
    xor g29980 ( n12725 , n28221 , n30740 );
    not g29981 ( n29847 , n10839 );
    or g29982 ( n10958 , n26884 , n15097 );
    xnor g29983 ( n16855 , n19778 , n1118 );
    or g29984 ( n31697 , n24061 , n14250 );
    nor g29985 ( n10743 , n23064 , n21377 );
    xnor g29986 ( n6596 , n28805 , n25960 );
    and g29987 ( n11593 , n9049 , n17987 );
    or g29988 ( n28128 , n2665 , n11950 );
    xnor g29989 ( n8455 , n170 , n19592 );
    xnor g29990 ( n1178 , n907 , n2258 );
    not g29991 ( n14104 , n30525 );
    nor g29992 ( n26942 , n20495 , n7209 );
    and g29993 ( n29865 , n3756 , n2310 );
    xnor g29994 ( n7881 , n23430 , n19524 );
    nor g29995 ( n23231 , n29705 , n28058 );
    or g29996 ( n15385 , n11258 , n17214 );
    not g29997 ( n5711 , n18518 );
    or g29998 ( n16013 , n13646 , n4738 );
    xnor g29999 ( n532 , n27153 , n9857 );
    or g30000 ( n4838 , n4551 , n28720 );
    or g30001 ( n30159 , n11629 , n967 );
    not g30002 ( n16369 , n30095 );
    not g30003 ( n27217 , n16963 );
    or g30004 ( n2505 , n5689 , n6576 );
    nor g30005 ( n6715 , n21124 , n15156 );
    or g30006 ( n22704 , n4214 , n9809 );
    xnor g30007 ( n2675 , n15396 , n12946 );
    xnor g30008 ( n16030 , n11648 , n18002 );
    or g30009 ( n1968 , n30118 , n3477 );
    and g30010 ( n26034 , n3604 , n2862 );
    buf g30011 ( n21310 , n27663 );
    or g30012 ( n14407 , n20568 , n10437 );
    not g30013 ( n28268 , n21231 );
    and g30014 ( n6649 , n21039 , n23342 );
    and g30015 ( n11334 , n15691 , n10621 );
    not g30016 ( n22596 , n30724 );
    or g30017 ( n23836 , n31091 , n26993 );
    not g30018 ( n11345 , n15436 );
    nor g30019 ( n17081 , n14100 , n9482 );
    xnor g30020 ( n1519 , n7823 , n24689 );
    not g30021 ( n15166 , n30394 );
    nor g30022 ( n7276 , n7316 , n16959 );
    not g30023 ( n17271 , n8415 );
    or g30024 ( n9169 , n350 , n14217 );
    or g30025 ( n14334 , n28240 , n31285 );
    or g30026 ( n21353 , n1634 , n940 );
    or g30027 ( n499 , n4494 , n15726 );
    xor g30028 ( n10928 , n2931 , n9592 );
    nor g30029 ( n21799 , n16308 , n29403 );
    or g30030 ( n16918 , n24029 , n11366 );
    and g30031 ( n4088 , n13068 , n7783 );
    and g30032 ( n9224 , n11484 , n26867 );
    not g30033 ( n4744 , n30405 );
    not g30034 ( n25209 , n1606 );
    not g30035 ( n17254 , n3195 );
    xnor g30036 ( n8067 , n12834 , n27757 );
    and g30037 ( n3607 , n15492 , n8285 );
    xnor g30038 ( n29692 , n29389 , n9620 );
    or g30039 ( n2194 , n16567 , n19016 );
    nor g30040 ( n21176 , n28058 , n20167 );
    or g30041 ( n27968 , n27763 , n10891 );
    xnor g30042 ( n6604 , n206 , n27022 );
    not g30043 ( n13507 , n5934 );
    nor g30044 ( n22006 , n11098 , n20067 );
    not g30045 ( n29955 , n3030 );
    nor g30046 ( n4417 , n3641 , n15684 );
    not g30047 ( n25296 , n4577 );
    xnor g30048 ( n29510 , n28506 , n30768 );
    xnor g30049 ( n20202 , n31303 , n12026 );
    not g30050 ( n20234 , n21346 );
    xnor g30051 ( n31566 , n14057 , n30850 );
    and g30052 ( n10106 , n25167 , n17917 );
    not g30053 ( n17628 , n1752 );
    not g30054 ( n3184 , n11736 );
    not g30055 ( n9033 , n3289 );
    xor g30056 ( n26657 , n11080 , n8042 );
    xnor g30057 ( n19762 , n11197 , n238 );
    or g30058 ( n26772 , n27920 , n4059 );
    or g30059 ( n6623 , n3076 , n7377 );
    or g30060 ( n9926 , n31113 , n18437 );
    xor g30061 ( n11981 , n26794 , n20181 );
    not g30062 ( n22691 , n21432 );
    xnor g30063 ( n27185 , n9627 , n30080 );
    not g30064 ( n3267 , n924 );
    not g30065 ( n15507 , n10507 );
    and g30066 ( n23132 , n12236 , n26815 );
    and g30067 ( n26357 , n1930 , n22482 );
    and g30068 ( n17113 , n24755 , n18738 );
    not g30069 ( n11502 , n28294 );
    not g30070 ( n20590 , n29998 );
    and g30071 ( n6879 , n30890 , n25290 );
    not g30072 ( n17319 , n26206 );
    or g30073 ( n21419 , n24184 , n15749 );
    not g30074 ( n15559 , n17149 );
    or g30075 ( n3612 , n28623 , n3264 );
    xor g30076 ( n12363 , n19995 , n8268 );
    not g30077 ( n26395 , n19538 );
    or g30078 ( n15959 , n18359 , n24642 );
    xnor g30079 ( n6507 , n3986 , n7014 );
    and g30080 ( n18195 , n18945 , n6108 );
    or g30081 ( n6693 , n30669 , n27321 );
    not g30082 ( n8285 , n30384 );
    not g30083 ( n12057 , n21141 );
    or g30084 ( n21779 , n16454 , n26389 );
    or g30085 ( n27812 , n7538 , n31939 );
    or g30086 ( n13094 , n26336 , n19479 );
    not g30087 ( n11870 , n3453 );
    nor g30088 ( n19349 , n20853 , n12567 );
    nor g30089 ( n26596 , n8924 , n21114 );
    or g30090 ( n6262 , n26686 , n15431 );
    not g30091 ( n13990 , n9693 );
    and g30092 ( n21967 , n14642 , n1263 );
    and g30093 ( n4338 , n7088 , n27228 );
    nor g30094 ( n26169 , n13968 , n15196 );
    or g30095 ( n15915 , n21656 , n19275 );
    and g30096 ( n24968 , n23766 , n17476 );
    not g30097 ( n31891 , n18955 );
    xnor g30098 ( n187 , n17352 , n7398 );
    or g30099 ( n25910 , n14086 , n27862 );
    not g30100 ( n2439 , n19375 );
    not g30101 ( n30465 , n24268 );
    nor g30102 ( n18363 , n27856 , n30714 );
    nor g30103 ( n2162 , n29717 , n19448 );
    not g30104 ( n23098 , n5719 );
    xnor g30105 ( n24774 , n26260 , n5218 );
    not g30106 ( n30271 , n28717 );
    not g30107 ( n16331 , n3297 );
    xnor g30108 ( n4988 , n29471 , n12668 );
    xnor g30109 ( n28558 , n3591 , n30769 );
    xnor g30110 ( n2673 , n20313 , n28983 );
    and g30111 ( n28221 , n21861 , n2351 );
    xnor g30112 ( n15512 , n14361 , n11905 );
    or g30113 ( n337 , n26870 , n26952 );
    not g30114 ( n10497 , n5642 );
    not g30115 ( n29679 , n11807 );
    or g30116 ( n17897 , n2835 , n20161 );
    not g30117 ( n27764 , n3596 );
    xnor g30118 ( n14515 , n15507 , n13348 );
    xnor g30119 ( n11457 , n3416 , n7026 );
    and g30120 ( n16327 , n14739 , n3027 );
    xnor g30121 ( n27572 , n7974 , n17398 );
    xnor g30122 ( n27508 , n26471 , n22846 );
    or g30123 ( n15910 , n24204 , n29622 );
    not g30124 ( n21613 , n7872 );
    and g30125 ( n13968 , n20891 , n2120 );
    xnor g30126 ( n22717 , n3520 , n25248 );
    not g30127 ( n9334 , n15550 );
    or g30128 ( n3045 , n15758 , n17843 );
    not g30129 ( n17437 , n22867 );
    or g30130 ( n21269 , n21085 , n8468 );
    or g30131 ( n29463 , n20442 , n20790 );
    or g30132 ( n1716 , n23209 , n9285 );
    or g30133 ( n26437 , n6387 , n913 );
    not g30134 ( n5770 , n757 );
    or g30135 ( n9261 , n25571 , n29814 );
    and g30136 ( n19511 , n25974 , n19133 );
    xnor g30137 ( n18939 , n28954 , n5883 );
    not g30138 ( n26091 , n734 );
    xnor g30139 ( n11148 , n14245 , n8053 );
    or g30140 ( n12833 , n20198 , n25525 );
    not g30141 ( n18848 , n3492 );
    and g30142 ( n23316 , n30653 , n26876 );
    not g30143 ( n6285 , n21047 );
    xnor g30144 ( n19557 , n19244 , n18877 );
    or g30145 ( n27726 , n5653 , n3103 );
    xnor g30146 ( n11649 , n26949 , n29467 );
    not g30147 ( n8839 , n26391 );
    or g30148 ( n12950 , n24605 , n18397 );
    or g30149 ( n27371 , n7204 , n6422 );
    xor g30150 ( n22968 , n1232 , n5128 );
    or g30151 ( n29244 , n9935 , n16804 );
    and g30152 ( n11656 , n5748 , n2499 );
    not g30153 ( n25541 , n13999 );
    not g30154 ( n11133 , n7594 );
    nor g30155 ( n27687 , n14373 , n3284 );
    not g30156 ( n24122 , n2199 );
    not g30157 ( n23801 , n4771 );
    not g30158 ( n26882 , n19891 );
    not g30159 ( n12351 , n11225 );
    xnor g30160 ( n25346 , n1157 , n2862 );
    xnor g30161 ( n4899 , n28792 , n9499 );
    nor g30162 ( n16195 , n8163 , n26371 );
    or g30163 ( n25138 , n20009 , n20072 );
    not g30164 ( n10980 , n2450 );
    not g30165 ( n13286 , n17863 );
    not g30166 ( n5556 , n30405 );
    not g30167 ( n9654 , n1048 );
    not g30168 ( n12602 , n19132 );
    and g30169 ( n9878 , n19175 , n23989 );
    not g30170 ( n14372 , n20629 );
    not g30171 ( n30928 , n19476 );
    or g30172 ( n10314 , n534 , n863 );
    or g30173 ( n17193 , n561 , n25265 );
    and g30174 ( n22015 , n31557 , n15405 );
    or g30175 ( n1462 , n13441 , n11693 );
    nor g30176 ( n1089 , n28562 , n11698 );
    not g30177 ( n3960 , n17580 );
    and g30178 ( n5582 , n20449 , n25061 );
    xnor g30179 ( n10965 , n16411 , n22316 );
    nor g30180 ( n11946 , n8827 , n30468 );
    not g30181 ( n14446 , n13356 );
    xnor g30182 ( n19980 , n22175 , n1882 );
    xnor g30183 ( n26233 , n6899 , n17375 );
    xnor g30184 ( n2451 , n30002 , n26894 );
    not g30185 ( n20642 , n4960 );
    not g30186 ( n15128 , n7641 );
    xnor g30187 ( n6041 , n29055 , n17302 );
    xnor g30188 ( n18251 , n8050 , n13959 );
    and g30189 ( n997 , n15239 , n1162 );
    xnor g30190 ( n7487 , n18566 , n24207 );
    or g30191 ( n16488 , n30339 , n11740 );
    not g30192 ( n17582 , n12078 );
    not g30193 ( n6972 , n7742 );
    xnor g30194 ( n24016 , n24919 , n811 );
    nor g30195 ( n26933 , n11666 , n9 );
    or g30196 ( n24364 , n22055 , n26288 );
    or g30197 ( n15932 , n12647 , n229 );
    and g30198 ( n10695 , n19906 , n605 );
    or g30199 ( n23269 , n23163 , n1832 );
    or g30200 ( n5364 , n13039 , n19541 );
    xnor g30201 ( n7942 , n20035 , n1202 );
    not g30202 ( n4140 , n19592 );
    not g30203 ( n20383 , n28068 );
    not g30204 ( n3278 , n23572 );
    and g30205 ( n6032 , n31312 , n31148 );
    or g30206 ( n18626 , n31094 , n28077 );
    nor g30207 ( n13146 , n11175 , n16385 );
    not g30208 ( n6607 , n4914 );
    xnor g30209 ( n2578 , n22094 , n21653 );
    xnor g30210 ( n20060 , n14484 , n5100 );
    and g30211 ( n21338 , n15701 , n38 );
    not g30212 ( n26658 , n23126 );
    nor g30213 ( n5629 , n13137 , n4539 );
    and g30214 ( n27834 , n25075 , n21666 );
    xnor g30215 ( n15471 , n15867 , n3895 );
    not g30216 ( n17519 , n10674 );
    and g30217 ( n9847 , n23698 , n28762 );
    not g30218 ( n21151 , n28034 );
    not g30219 ( n19445 , n10630 );
    or g30220 ( n16251 , n12014 , n30392 );
    and g30221 ( n21753 , n6877 , n3811 );
    and g30222 ( n9014 , n31843 , n16933 );
    and g30223 ( n11993 , n5472 , n16756 );
    not g30224 ( n13922 , n9725 );
    not g30225 ( n2779 , n3515 );
    or g30226 ( n23168 , n4527 , n25463 );
    not g30227 ( n9816 , n17286 );
    xnor g30228 ( n30163 , n30054 , n20978 );
    or g30229 ( n20457 , n6980 , n20011 );
    or g30230 ( n31834 , n26594 , n15961 );
    xnor g30231 ( n1281 , n9268 , n5499 );
    and g30232 ( n31683 , n17936 , n22655 );
    not g30233 ( n26993 , n20453 );
    or g30234 ( n4679 , n25603 , n18169 );
    or g30235 ( n26316 , n238 , n22112 );
    not g30236 ( n27637 , n3326 );
    not g30237 ( n5067 , n23074 );
    not g30238 ( n7608 , n31798 );
    not g30239 ( n26500 , n5455 );
    or g30240 ( n3380 , n23231 , n789 );
    xnor g30241 ( n22751 , n7414 , n8584 );
    xnor g30242 ( n452 , n10788 , n30896 );
    or g30243 ( n7918 , n21852 , n164 );
    not g30244 ( n8124 , n30794 );
    or g30245 ( n155 , n2189 , n2622 );
    xnor g30246 ( n18444 , n12790 , n21472 );
    and g30247 ( n22071 , n26618 , n9919 );
    nor g30248 ( n17425 , n24199 , n23687 );
    xnor g30249 ( n22433 , n25276 , n14967 );
    xnor g30250 ( n21445 , n30549 , n6874 );
    and g30251 ( n17626 , n16768 , n3016 );
    and g30252 ( n30035 , n25271 , n11154 );
    not g30253 ( n29272 , n3971 );
    or g30254 ( n17351 , n18653 , n4690 );
    not g30255 ( n31178 , n26585 );
    and g30256 ( n3103 , n6004 , n17120 );
    xor g30257 ( n12122 , n231 , n6651 );
    or g30258 ( n13390 , n8642 , n16838 );
    or g30259 ( n24690 , n12186 , n25715 );
    or g30260 ( n805 , n23300 , n11988 );
    xnor g30261 ( n29049 , n17617 , n6603 );
    xnor g30262 ( n7650 , n29523 , n19933 );
    and g30263 ( n25274 , n29936 , n4054 );
    not g30264 ( n12146 , n21436 );
    xnor g30265 ( n23956 , n19726 , n24848 );
    xnor g30266 ( n4562 , n23541 , n1635 );
    and g30267 ( n450 , n4801 , n5843 );
    or g30268 ( n1287 , n14493 , n5239 );
    xor g30269 ( n31325 , n6984 , n4082 );
    and g30270 ( n26452 , n6605 , n1253 );
    and g30271 ( n16828 , n12847 , n29598 );
    nor g30272 ( n17764 , n21496 , n14843 );
    and g30273 ( n9007 , n21380 , n28964 );
    xnor g30274 ( n10959 , n26749 , n30287 );
    xor g30275 ( n3069 , n9907 , n24083 );
    nor g30276 ( n31367 , n30934 , n17437 );
    or g30277 ( n4580 , n2331 , n24181 );
    not g30278 ( n5506 , n31327 );
    or g30279 ( n4505 , n25238 , n1356 );
    not g30280 ( n9070 , n28934 );
    and g30281 ( n5789 , n28055 , n21508 );
    and g30282 ( n12581 , n31796 , n13769 );
    not g30283 ( n19157 , n7109 );
    and g30284 ( n13342 , n1286 , n20999 );
    or g30285 ( n25542 , n15496 , n8374 );
    nor g30286 ( n30825 , n27455 , n21879 );
    xnor g30287 ( n27223 , n6638 , n15509 );
    or g30288 ( n7612 , n30173 , n31640 );
    or g30289 ( n30671 , n25647 , n11151 );
    and g30290 ( n31673 , n5634 , n28620 );
    xnor g30291 ( n22100 , n28154 , n8987 );
    not g30292 ( n30434 , n24131 );
    not g30293 ( n14805 , n3946 );
    not g30294 ( n9137 , n3688 );
    or g30295 ( n8294 , n10485 , n15550 );
    and g30296 ( n24671 , n5294 , n6145 );
    not g30297 ( n24274 , n9168 );
    not g30298 ( n23183 , n27910 );
    and g30299 ( n20152 , n17958 , n22190 );
    xnor g30300 ( n17601 , n21662 , n22302 );
    xnor g30301 ( n24185 , n133 , n6768 );
    xnor g30302 ( n30153 , n26402 , n18128 );
    buf g30303 ( n20156 , n10067 );
    not g30304 ( n27901 , n27917 );
    xnor g30305 ( n5934 , n20586 , n20089 );
    xnor g30306 ( n30579 , n6068 , n4393 );
    or g30307 ( n19126 , n27390 , n23129 );
    not g30308 ( n6342 , n28213 );
    nor g30309 ( n9000 , n23207 , n11215 );
    and g30310 ( n31578 , n18385 , n31725 );
    buf g30311 ( n12857 , n17596 );
    or g30312 ( n23318 , n15530 , n29431 );
    xnor g30313 ( n29649 , n1099 , n21414 );
    nor g30314 ( n23027 , n16061 , n29539 );
    xnor g30315 ( n23538 , n19288 , n963 );
    nor g30316 ( n11147 , n25461 , n17135 );
    xnor g30317 ( n13364 , n7373 , n8787 );
    xnor g30318 ( n6206 , n7563 , n757 );
    not g30319 ( n22976 , n16409 );
    or g30320 ( n39 , n19347 , n13645 );
    xnor g30321 ( n16481 , n20984 , n19 );
    xor g30322 ( n22787 , n24787 , n998 );
    or g30323 ( n16136 , n20565 , n10563 );
    xnor g30324 ( n15194 , n17349 , n36 );
    not g30325 ( n28132 , n32025 );
    not g30326 ( n21079 , n18651 );
    not g30327 ( n7934 , n5299 );
    and g30328 ( n19874 , n24039 , n10890 );
    not g30329 ( n29015 , n1687 );
    xnor g30330 ( n29248 , n31977 , n17163 );
    nor g30331 ( n19482 , n757 , n26659 );
    not g30332 ( n13157 , n14796 );
    and g30333 ( n135 , n10191 , n29258 );
    not g30334 ( n470 , n15211 );
    xnor g30335 ( n26227 , n456 , n28825 );
    or g30336 ( n17231 , n24088 , n12626 );
    or g30337 ( n22984 , n27790 , n26110 );
    not g30338 ( n4595 , n20797 );
    or g30339 ( n18456 , n8950 , n7724 );
    not g30340 ( n12674 , n22411 );
    nor g30341 ( n5618 , n10237 , n28247 );
    not g30342 ( n2116 , n19211 );
    not g30343 ( n8778 , n12338 );
    not g30344 ( n6006 , n22903 );
    or g30345 ( n11546 , n11133 , n21773 );
    xnor g30346 ( n7464 , n27910 , n1783 );
    not g30347 ( n31954 , n24724 );
    or g30348 ( n22195 , n23157 , n10807 );
    and g30349 ( n692 , n21115 , n1845 );
    not g30350 ( n12042 , n20743 );
    not g30351 ( n17357 , n23293 );
    xnor g30352 ( n28085 , n13582 , n4384 );
    xnor g30353 ( n5396 , n29280 , n29117 );
    or g30354 ( n5139 , n2498 , n21587 );
    not g30355 ( n63 , n15413 );
    and g30356 ( n14791 , n6384 , n30227 );
    not g30357 ( n28635 , n28998 );
    xnor g30358 ( n22979 , n27188 , n27157 );
    xnor g30359 ( n2407 , n17884 , n27077 );
    not g30360 ( n10848 , n2450 );
    and g30361 ( n4638 , n955 , n25632 );
    and g30362 ( n902 , n25025 , n25959 );
    or g30363 ( n4627 , n27161 , n32034 );
    or g30364 ( n18217 , n22762 , n30518 );
    and g30365 ( n24925 , n30662 , n11731 );
    xnor g30366 ( n20097 , n25089 , n8988 );
    not g30367 ( n18763 , n6492 );
    not g30368 ( n6804 , n21465 );
    or g30369 ( n19722 , n5200 , n30721 );
    not g30370 ( n7656 , n28953 );
    and g30371 ( n24855 , n6557 , n21498 );
    or g30372 ( n1778 , n8994 , n12522 );
    xnor g30373 ( n26653 , n8390 , n6437 );
    not g30374 ( n12604 , n24908 );
    and g30375 ( n15098 , n24479 , n5406 );
    xnor g30376 ( n26980 , n10154 , n29559 );
    or g30377 ( n560 , n7241 , n19572 );
    xnor g30378 ( n28745 , n19720 , n10034 );
    xnor g30379 ( n13748 , n4257 , n11262 );
    or g30380 ( n4452 , n1842 , n25277 );
    and g30381 ( n15150 , n15443 , n2003 );
    or g30382 ( n9132 , n15769 , n11191 );
    or g30383 ( n23321 , n9509 , n16713 );
    or g30384 ( n27588 , n26950 , n13531 );
    and g30385 ( n6627 , n16041 , n27069 );
    or g30386 ( n16046 , n12274 , n12149 );
    xnor g30387 ( n10922 , n8343 , n31319 );
    nor g30388 ( n28879 , n26029 , n26963 );
    and g30389 ( n18694 , n8937 , n670 );
    xnor g30390 ( n23013 , n29248 , n20655 );
    xnor g30391 ( n30982 , n10510 , n26780 );
    and g30392 ( n17744 , n5821 , n23244 );
    or g30393 ( n18228 , n27457 , n6786 );
    and g30394 ( n28025 , n26609 , n21186 );
    and g30395 ( n7410 , n26572 , n20706 );
    or g30396 ( n30749 , n25388 , n21399 );
    nor g30397 ( n10458 , n23552 , n251 );
    xnor g30398 ( n30186 , n23717 , n19385 );
    not g30399 ( n30247 , n12009 );
    nor g30400 ( n15034 , n13151 , n13799 );
    xor g30401 ( n7894 , n4760 , n21771 );
    not g30402 ( n30468 , n18447 );
    and g30403 ( n10499 , n29827 , n31027 );
    and g30404 ( n23290 , n2538 , n31146 );
    xnor g30405 ( n28836 , n13062 , n1346 );
    or g30406 ( n15451 , n27709 , n3954 );
    xor g30407 ( n24515 , n27006 , n18445 );
    not g30408 ( n9371 , n4445 );
    xnor g30409 ( n28808 , n22579 , n17227 );
    not g30410 ( n26183 , n23405 );
    or g30411 ( n4976 , n6167 , n20147 );
    not g30412 ( n23659 , n3614 );
    not g30413 ( n4033 , n1796 );
    not g30414 ( n31460 , n10148 );
    not g30415 ( n28610 , n29293 );
    not g30416 ( n19737 , n3265 );
    and g30417 ( n24290 , n5188 , n28735 );
    and g30418 ( n9913 , n28074 , n22621 );
    or g30419 ( n29302 , n28875 , n18881 );
    or g30420 ( n15919 , n909 , n27382 );
    not g30421 ( n7141 , n16654 );
    not g30422 ( n18842 , n20822 );
    or g30423 ( n23570 , n15374 , n11932 );
    and g30424 ( n21532 , n5807 , n26411 );
    xnor g30425 ( n2146 , n20581 , n23309 );
    nor g30426 ( n12905 , n2444 , n21186 );
    or g30427 ( n10401 , n24679 , n28129 );
    not g30428 ( n30461 , n6371 );
    or g30429 ( n23233 , n22449 , n28575 );
    xnor g30430 ( n2476 , n5792 , n9321 );
    or g30431 ( n16547 , n17543 , n12081 );
    and g30432 ( n478 , n4151 , n17718 );
    not g30433 ( n15315 , n1787 );
    or g30434 ( n1757 , n10419 , n26835 );
    not g30435 ( n5041 , n17894 );
    xnor g30436 ( n1031 , n20073 , n31619 );
    xor g30437 ( n12936 , n22521 , n14792 );
    not g30438 ( n16867 , n27207 );
    xnor g30439 ( n8847 , n26793 , n23097 );
    not g30440 ( n6984 , n27322 );
    xnor g30441 ( n31361 , n23803 , n10649 );
    and g30442 ( n3089 , n7853 , n24243 );
    or g30443 ( n30086 , n14871 , n15490 );
    xnor g30444 ( n19584 , n13191 , n30971 );
    or g30445 ( n23952 , n3472 , n7629 );
    not g30446 ( n17561 , n8714 );
    or g30447 ( n4308 , n3996 , n3485 );
    or g30448 ( n17311 , n22373 , n4319 );
    nor g30449 ( n30265 , n25488 , n2753 );
    nor g30450 ( n16422 , n11306 , n20579 );
    not g30451 ( n9343 , n7215 );
    not g30452 ( n1751 , n27168 );
    and g30453 ( n12156 , n13692 , n19636 );
    not g30454 ( n2385 , n23339 );
    xnor g30455 ( n29314 , n22320 , n13154 );
    or g30456 ( n176 , n25608 , n7161 );
    xnor g30457 ( n30156 , n3597 , n6745 );
    and g30458 ( n14369 , n18780 , n10430 );
    nor g30459 ( n22628 , n11400 , n31752 );
    or g30460 ( n28823 , n11563 , n17575 );
    and g30461 ( n15909 , n1012 , n30669 );
    nor g30462 ( n26612 , n30045 , n6422 );
    xnor g30463 ( n2700 , n3243 , n28475 );
    nor g30464 ( n2635 , n22927 , n13136 );
    xnor g30465 ( n12256 , n18900 , n20116 );
    xnor g30466 ( n1024 , n7072 , n25714 );
    xnor g30467 ( n4709 , n5854 , n26052 );
    not g30468 ( n18866 , n28870 );
    xnor g30469 ( n1220 , n20915 , n20074 );
    xnor g30470 ( n1646 , n7446 , n29304 );
    not g30471 ( n31276 , n12130 );
    not g30472 ( n22088 , n6168 );
    and g30473 ( n8472 , n23671 , n8640 );
    xnor g30474 ( n3839 , n5384 , n2483 );
    and g30475 ( n20762 , n11790 , n11125 );
    or g30476 ( n19250 , n10349 , n31213 );
    xnor g30477 ( n980 , n30237 , n22696 );
    not g30478 ( n30557 , n25245 );
    not g30479 ( n2722 , n21670 );
    not g30480 ( n19440 , n17713 );
    or g30481 ( n7973 , n25605 , n1056 );
    or g30482 ( n27499 , n12679 , n25604 );
    xnor g30483 ( n29795 , n23003 , n18300 );
    xnor g30484 ( n16203 , n12067 , n17763 );
    and g30485 ( n12542 , n1386 , n17811 );
    xnor g30486 ( n30063 , n31561 , n28447 );
    xnor g30487 ( n9633 , n11554 , n4358 );
    nor g30488 ( n3679 , n12072 , n18534 );
    xnor g30489 ( n26542 , n10488 , n12688 );
    or g30490 ( n19895 , n30149 , n2201 );
    not g30491 ( n11979 , n7138 );
    or g30492 ( n27245 , n24711 , n30098 );
    xnor g30493 ( n24398 , n12005 , n2530 );
    or g30494 ( n1135 , n6874 , n30549 );
    and g30495 ( n31253 , n8979 , n12311 );
    not g30496 ( n15258 , n25774 );
    not g30497 ( n21293 , n11215 );
    nor g30498 ( n12521 , n24911 , n14057 );
    nor g30499 ( n4001 , n9145 , n25532 );
    xnor g30500 ( n16594 , n18203 , n13859 );
    or g30501 ( n5324 , n11360 , n20412 );
    or g30502 ( n18422 , n21100 , n31816 );
    or g30503 ( n31908 , n24023 , n4372 );
    or g30504 ( n23766 , n27118 , n3279 );
    and g30505 ( n16505 , n15314 , n25439 );
    and g30506 ( n25650 , n21710 , n24383 );
    xnor g30507 ( n25714 , n1736 , n15272 );
    xnor g30508 ( n6386 , n4718 , n10055 );
    not g30509 ( n4525 , n14711 );
    xnor g30510 ( n7884 , n18081 , n23858 );
    nor g30511 ( n1216 , n13065 , n17951 );
    or g30512 ( n20266 , n21186 , n26609 );
    xnor g30513 ( n23806 , n13307 , n4663 );
    or g30514 ( n24658 , n21999 , n8543 );
    not g30515 ( n4696 , n21302 );
    or g30516 ( n378 , n22877 , n1981 );
    xnor g30517 ( n11394 , n11144 , n16290 );
    not g30518 ( n25628 , n31411 );
    and g30519 ( n11150 , n18016 , n8481 );
    not g30520 ( n13267 , n6027 );
    xnor g30521 ( n14418 , n377 , n24093 );
    not g30522 ( n14335 , n23522 );
    and g30523 ( n25941 , n11310 , n1578 );
    and g30524 ( n16326 , n6725 , n1366 );
    xnor g30525 ( n20894 , n25307 , n21187 );
    nor g30526 ( n28727 , n6864 , n18689 );
    xnor g30527 ( n20827 , n13195 , n19856 );
    not g30528 ( n23503 , n474 );
    or g30529 ( n21145 , n14968 , n18563 );
    xnor g30530 ( n5753 , n9989 , n4972 );
    not g30531 ( n31102 , n30830 );
    and g30532 ( n13178 , n18459 , n26638 );
    xnor g30533 ( n18728 , n23960 , n28081 );
    and g30534 ( n29281 , n1183 , n21482 );
    or g30535 ( n23106 , n11703 , n4066 );
    and g30536 ( n18250 , n16834 , n9283 );
    and g30537 ( n16923 , n3126 , n26692 );
    xnor g30538 ( n13504 , n22676 , n28598 );
    xnor g30539 ( n26919 , n11890 , n2389 );
    or g30540 ( n8629 , n6552 , n29540 );
    xnor g30541 ( n27872 , n12701 , n25121 );
    nor g30542 ( n18949 , n6957 , n28258 );
    xnor g30543 ( n125 , n18594 , n20316 );
    and g30544 ( n6781 , n16751 , n31003 );
    not g30545 ( n10905 , n11289 );
    xnor g30546 ( n15482 , n18496 , n16558 );
    and g30547 ( n19381 , n29459 , n20331 );
    or g30548 ( n17999 , n30711 , n5491 );
    or g30549 ( n25712 , n29375 , n18954 );
    and g30550 ( n23121 , n20488 , n23941 );
    xnor g30551 ( n26213 , n19353 , n8841 );
    or g30552 ( n15515 , n29111 , n29026 );
    xnor g30553 ( n4148 , n26894 , n6874 );
    xnor g30554 ( n11841 , n13927 , n23400 );
    not g30555 ( n19887 , n20510 );
    nor g30556 ( n25098 , n6331 , n8321 );
    not g30557 ( n27067 , n812 );
    xnor g30558 ( n12556 , n23261 , n2994 );
    buf g30559 ( n6750 , n6659 );
    and g30560 ( n14213 , n5258 , n19108 );
    not g30561 ( n6472 , n25276 );
    nor g30562 ( n6387 , n18645 , n18850 );
    or g30563 ( n22179 , n27814 , n19005 );
    xnor g30564 ( n25627 , n19091 , n28562 );
    xnor g30565 ( n21217 , n21494 , n31783 );
    xnor g30566 ( n8609 , n18522 , n3905 );
    xnor g30567 ( n3962 , n15962 , n19790 );
    or g30568 ( n17970 , n13210 , n9663 );
    or g30569 ( n16394 , n20690 , n17953 );
    not g30570 ( n15348 , n30458 );
    xnor g30571 ( n31864 , n21905 , n7674 );
    and g30572 ( n24853 , n1543 , n26598 );
    and g30573 ( n6742 , n1454 , n21371 );
    and g30574 ( n4669 , n2522 , n23611 );
    not g30575 ( n3745 , n21561 );
    xnor g30576 ( n26576 , n15356 , n30162 );
    or g30577 ( n30871 , n15588 , n6009 );
    or g30578 ( n21859 , n13144 , n3504 );
    not g30579 ( n20599 , n25208 );
    not g30580 ( n13022 , n29617 );
    xnor g30581 ( n14368 , n19708 , n30065 );
    xnor g30582 ( n10684 , n29449 , n2502 );
    xnor g30583 ( n29051 , n2354 , n15358 );
    xnor g30584 ( n16563 , n13099 , n26123 );
    or g30585 ( n24646 , n17182 , n7750 );
    xnor g30586 ( n19676 , n14830 , n1432 );
    or g30587 ( n22048 , n28417 , n11341 );
    xnor g30588 ( n1999 , n15541 , n29640 );
    not g30589 ( n20216 , n16281 );
    or g30590 ( n16952 , n10955 , n14070 );
    or g30591 ( n16628 , n18976 , n6855 );
    or g30592 ( n12382 , n30155 , n31909 );
    nor g30593 ( n11548 , n17019 , n16914 );
    or g30594 ( n24502 , n11564 , n11751 );
    or g30595 ( n20375 , n30004 , n31953 );
    and g30596 ( n6222 , n8780 , n25846 );
    or g30597 ( n2269 , n3856 , n984 );
    and g30598 ( n9644 , n12555 , n26427 );
    xnor g30599 ( n27310 , n16113 , n23115 );
    xnor g30600 ( n4396 , n10880 , n11584 );
    not g30601 ( n10220 , n16607 );
    xor g30602 ( n4187 , n25874 , n11180 );
    and g30603 ( n28429 , n1584 , n21117 );
    and g30604 ( n24719 , n23028 , n15316 );
    xnor g30605 ( n27488 , n9770 , n20977 );
    not g30606 ( n12865 , n17025 );
    xnor g30607 ( n26415 , n6877 , n7833 );
    xor g30608 ( n28909 , n22339 , n24449 );
    not g30609 ( n31671 , n16871 );
    and g30610 ( n7874 , n9950 , n29074 );
    or g30611 ( n14866 , n21146 , n6081 );
    and g30612 ( n28011 , n23819 , n1146 );
    not g30613 ( n7084 , n27083 );
    and g30614 ( n9836 , n28234 , n17851 );
    or g30615 ( n7989 , n20486 , n13519 );
    and g30616 ( n17282 , n12466 , n8146 );
    not g30617 ( n17069 , n4220 );
    xnor g30618 ( n29842 , n14223 , n25661 );
    not g30619 ( n16492 , n1039 );
    and g30620 ( n20958 , n29560 , n23026 );
    xor g30621 ( n9854 , n19824 , n10299 );
    and g30622 ( n6832 , n9108 , n1809 );
    or g30623 ( n17107 , n27687 , n11578 );
    not g30624 ( n30686 , n12146 );
    and g30625 ( n6109 , n7361 , n13522 );
    not g30626 ( n21668 , n7129 );
    or g30627 ( n15428 , n23134 , n2247 );
    not g30628 ( n7644 , n21800 );
    xnor g30629 ( n28579 , n11117 , n9209 );
    and g30630 ( n8530 , n26221 , n30517 );
    not g30631 ( n15793 , n30685 );
    not g30632 ( n8978 , n29756 );
    nor g30633 ( n17733 , n27373 , n499 );
    and g30634 ( n13633 , n12281 , n19551 );
    not g30635 ( n17729 , n29285 );
    not g30636 ( n11139 , n859 );
    xnor g30637 ( n18292 , n10992 , n22695 );
    not g30638 ( n11093 , n797 );
    xnor g30639 ( n6392 , n112 , n5575 );
    xnor g30640 ( n4743 , n5363 , n26891 );
    or g30641 ( n22267 , n26745 , n18197 );
    not g30642 ( n4637 , n22442 );
    not g30643 ( n27701 , n20870 );
    or g30644 ( n5093 , n28504 , n7174 );
    not g30645 ( n28294 , n8312 );
    not g30646 ( n31664 , n14121 );
    or g30647 ( n4713 , n31633 , n23944 );
    xnor g30648 ( n11560 , n4157 , n30587 );
    and g30649 ( n20025 , n3691 , n30514 );
    or g30650 ( n15023 , n25059 , n10726 );
    nor g30651 ( n31580 , n10589 , n30893 );
    or g30652 ( n19227 , n473 , n10260 );
    xnor g30653 ( n19919 , n18478 , n18090 );
    or g30654 ( n7450 , n14954 , n17145 );
    nor g30655 ( n5611 , n11611 , n4227 );
    not g30656 ( n14757 , n17317 );
    not g30657 ( n20821 , n26217 );
    not g30658 ( n18833 , n3306 );
    not g30659 ( n19155 , n30401 );
    xnor g30660 ( n31020 , n23109 , n15619 );
    xnor g30661 ( n1845 , n13627 , n29595 );
    and g30662 ( n31087 , n8169 , n20083 );
    nor g30663 ( n26622 , n19505 , n22142 );
    not g30664 ( n9895 , n18543 );
    not g30665 ( n27208 , n9070 );
    and g30666 ( n1019 , n13624 , n1295 );
    not g30667 ( n3616 , n19113 );
    xor g30668 ( n24876 , n6081 , n21689 );
    or g30669 ( n12977 , n19218 , n26376 );
    not g30670 ( n26060 , n19590 );
    not g30671 ( n28111 , n20279 );
    and g30672 ( n30355 , n23509 , n18304 );
    nor g30673 ( n9287 , n21824 , n8722 );
    xnor g30674 ( n152 , n26480 , n17751 );
    not g30675 ( n2446 , n6135 );
    xnor g30676 ( n6917 , n8720 , n12803 );
    xnor g30677 ( n24262 , n29896 , n7641 );
    and g30678 ( n27686 , n9162 , n15936 );
    or g30679 ( n30073 , n2583 , n6769 );
    not g30680 ( n26607 , n26541 );
    xnor g30681 ( n8217 , n554 , n23232 );
    and g30682 ( n816 , n22720 , n12413 );
    not g30683 ( n7915 , n31906 );
    xnor g30684 ( n13572 , n15495 , n17368 );
    not g30685 ( n2196 , n7200 );
    nor g30686 ( n6948 , n20236 , n23518 );
    and g30687 ( n9024 , n21130 , n1091 );
    not g30688 ( n21291 , n22835 );
    not g30689 ( n4031 , n18318 );
    xnor g30690 ( n27410 , n27852 , n27029 );
    and g30691 ( n12040 , n15267 , n27819 );
    not g30692 ( n11928 , n14894 );
    and g30693 ( n24778 , n21247 , n12736 );
    nor g30694 ( n308 , n15756 , n9371 );
    not g30695 ( n9061 , n16006 );
    xnor g30696 ( n28815 , n1271 , n24115 );
    or g30697 ( n9725 , n23518 , n16213 );
    nor g30698 ( n9595 , n31828 , n17370 );
    xnor g30699 ( n16861 , n13873 , n29806 );
    not g30700 ( n29436 , n30728 );
    nor g30701 ( n21317 , n2869 , n1652 );
    xnor g30702 ( n16361 , n20610 , n5673 );
    and g30703 ( n1158 , n18618 , n4333 );
    not g30704 ( n18498 , n2317 );
    not g30705 ( n20756 , n17100 );
    nor g30706 ( n15168 , n17310 , n10041 );
    nor g30707 ( n12328 , n12390 , n15764 );
    xnor g30708 ( n151 , n4897 , n16685 );
    nor g30709 ( n11182 , n12312 , n3787 );
    or g30710 ( n23219 , n2148 , n2374 );
    nor g30711 ( n25094 , n10477 , n956 );
    or g30712 ( n23329 , n8068 , n1289 );
    not g30713 ( n18789 , n8936 );
    xnor g30714 ( n20767 , n14954 , n22665 );
    or g30715 ( n2909 , n29132 , n9561 );
    or g30716 ( n13522 , n11984 , n3367 );
    not g30717 ( n6842 , n22375 );
    not g30718 ( n3818 , n4907 );
    and g30719 ( n25733 , n9829 , n17302 );
    xnor g30720 ( n17439 , n21792 , n28168 );
    not g30721 ( n25874 , n3810 );
    or g30722 ( n955 , n11779 , n31687 );
    and g30723 ( n21856 , n24501 , n11515 );
    or g30724 ( n22932 , n4054 , n29936 );
    not g30725 ( n8576 , n11065 );
    not g30726 ( n15390 , n20291 );
    and g30727 ( n19347 , n28930 , n23469 );
    not g30728 ( n4768 , n19236 );
    xor g30729 ( n11804 , n12469 , n28517 );
    xnor g30730 ( n23136 , n5413 , n31215 );
    or g30731 ( n23000 , n13043 , n12809 );
    or g30732 ( n6185 , n1473 , n22946 );
    not g30733 ( n22560 , n6010 );
    and g30734 ( n11146 , n23329 , n11754 );
    or g30735 ( n6158 , n20400 , n27997 );
    not g30736 ( n29028 , n12371 );
    not g30737 ( n25896 , n9831 );
    or g30738 ( n27329 , n13991 , n25964 );
    not g30739 ( n257 , n18389 );
    xnor g30740 ( n25976 , n10100 , n13018 );
    not g30741 ( n7514 , n256 );
    or g30742 ( n10225 , n4793 , n12507 );
    or g30743 ( n22847 , n5027 , n27270 );
    xnor g30744 ( n20522 , n15178 , n3641 );
    xnor g30745 ( n30373 , n22282 , n23925 );
    and g30746 ( n31487 , n3903 , n11982 );
    and g30747 ( n13606 , n16469 , n7250 );
    xnor g30748 ( n18773 , n20663 , n16660 );
    and g30749 ( n20258 , n3666 , n15982 );
    xnor g30750 ( n22466 , n25391 , n8619 );
    xnor g30751 ( n27904 , n26826 , n13764 );
    nor g30752 ( n16089 , n16970 , n27136 );
    or g30753 ( n2197 , n7533 , n12510 );
    or g30754 ( n24303 , n22824 , n13915 );
    nor g30755 ( n20887 , n13220 , n29384 );
    or g30756 ( n15217 , n28515 , n20783 );
    and g30757 ( n21560 , n17314 , n2972 );
    and g30758 ( n16913 , n5875 , n27283 );
    not g30759 ( n30346 , n5238 );
    or g30760 ( n3807 , n1204 , n22345 );
    xnor g30761 ( n15240 , n15392 , n29890 );
    not g30762 ( n18566 , n1812 );
    and g30763 ( n9114 , n9815 , n24106 );
    xnor g30764 ( n15053 , n8954 , n9705 );
    and g30765 ( n19189 , n28949 , n21183 );
    not g30766 ( n6871 , n6534 );
    not g30767 ( n21245 , n24918 );
    nor g30768 ( n6773 , n6882 , n8800 );
    not g30769 ( n24423 , n31330 );
    nor g30770 ( n7895 , n3447 , n28979 );
    or g30771 ( n12608 , n29284 , n24547 );
    not g30772 ( n22011 , n13130 );
    not g30773 ( n7592 , n16783 );
    xor g30774 ( n30549 , n12098 , n3106 );
    or g30775 ( n24952 , n18253 , n2510 );
    or g30776 ( n12956 , n31090 , n6350 );
    xnor g30777 ( n18252 , n30865 , n6295 );
    not g30778 ( n19254 , n11425 );
    not g30779 ( n7897 , n13142 );
    nor g30780 ( n11473 , n12496 , n23029 );
    or g30781 ( n11895 , n12712 , n30608 );
    not g30782 ( n24241 , n31695 );
    xnor g30783 ( n19080 , n31308 , n2420 );
    or g30784 ( n29381 , n11548 , n16969 );
    xnor g30785 ( n3282 , n12006 , n6537 );
    xnor g30786 ( n13976 , n14642 , n11915 );
    or g30787 ( n6203 , n3883 , n20086 );
    and g30788 ( n31730 , n11289 , n15009 );
    and g30789 ( n31308 , n3779 , n26679 );
    xnor g30790 ( n13963 , n4014 , n3333 );
    not g30791 ( n10528 , n5812 );
    not g30792 ( n22041 , n714 );
    or g30793 ( n24533 , n9613 , n19496 );
    and g30794 ( n15218 , n14151 , n30041 );
    not g30795 ( n14696 , n28121 );
    not g30796 ( n21227 , n12111 );
    xnor g30797 ( n13293 , n16094 , n22935 );
    xnor g30798 ( n2275 , n31914 , n27538 );
    not g30799 ( n8542 , n21080 );
    nor g30800 ( n19192 , n31035 , n53 );
    or g30801 ( n383 , n14363 , n12605 );
    xnor g30802 ( n12467 , n23504 , n30838 );
    not g30803 ( n22392 , n7064 );
    xnor g30804 ( n11701 , n28723 , n16156 );
    or g30805 ( n22297 , n27927 , n12097 );
    or g30806 ( n2566 , n30936 , n1698 );
    and g30807 ( n12059 , n4775 , n17175 );
    or g30808 ( n15956 , n13690 , n22349 );
    not g30809 ( n8722 , n2963 );
    or g30810 ( n12247 , n31426 , n5187 );
    not g30811 ( n12519 , n30161 );
    and g30812 ( n13323 , n13857 , n2704 );
    and g30813 ( n29735 , n19709 , n23924 );
    not g30814 ( n1534 , n18750 );
    or g30815 ( n18223 , n12777 , n1859 );
    or g30816 ( n27825 , n15201 , n1910 );
    or g30817 ( n14285 , n20657 , n31007 );
    or g30818 ( n5585 , n25413 , n6160 );
    xnor g30819 ( n4215 , n18815 , n6784 );
    not g30820 ( n20961 , n4023 );
    or g30821 ( n12289 , n3599 , n13331 );
    and g30822 ( n17887 , n27457 , n11502 );
    nor g30823 ( n846 , n9011 , n21186 );
    xnor g30824 ( n15603 , n3422 , n10847 );
    or g30825 ( n7100 , n11261 , n3099 );
    and g30826 ( n7629 , n22769 , n8886 );
    not g30827 ( n18119 , n12672 );
    and g30828 ( n11623 , n22604 , n14476 );
    or g30829 ( n17606 , n24534 , n15899 );
    not g30830 ( n14964 , n16649 );
    and g30831 ( n22153 , n14027 , n5342 );
    xnor g30832 ( n13601 , n19282 , n28402 );
    and g30833 ( n28430 , n18505 , n1409 );
    or g30834 ( n14384 , n27608 , n20123 );
    or g30835 ( n12586 , n26852 , n31315 );
    or g30836 ( n4043 , n1723 , n11830 );
    xnor g30837 ( n16529 , n508 , n27591 );
    xnor g30838 ( n12374 , n25471 , n31368 );
    and g30839 ( n23066 , n28229 , n2318 );
    not g30840 ( n3322 , n8531 );
    or g30841 ( n20963 , n397 , n30453 );
    or g30842 ( n17301 , n18207 , n27491 );
    not g30843 ( n12342 , n7362 );
    not g30844 ( n28831 , n3978 );
    or g30845 ( n6605 , n8504 , n22439 );
    xnor g30846 ( n24860 , n2856 , n969 );
    not g30847 ( n24867 , n19988 );
    not g30848 ( n14649 , n1131 );
    xnor g30849 ( n9291 , n10627 , n8260 );
    xnor g30850 ( n565 , n17642 , n21135 );
    xnor g30851 ( n27023 , n8644 , n10380 );
    not g30852 ( n14280 , n1002 );
    xnor g30853 ( n23443 , n8014 , n107 );
    and g30854 ( n13466 , n22293 , n15913 );
    and g30855 ( n20628 , n9547 , n4346 );
    xor g30856 ( n27975 , n11203 , n22665 );
    or g30857 ( n20179 , n12313 , n20945 );
    and g30858 ( n11580 , n9498 , n14670 );
    xnor g30859 ( n13923 , n5360 , n27034 );
    not g30860 ( n498 , n18310 );
    nor g30861 ( n20049 , n18836 , n22870 );
    not g30862 ( n7270 , n29363 );
    or g30863 ( n8533 , n1493 , n24855 );
    nor g30864 ( n18093 , n12711 , n17355 );
    and g30865 ( n28364 , n16879 , n31295 );
    not g30866 ( n9852 , n2677 );
    xnor g30867 ( n26565 , n25203 , n7983 );
    and g30868 ( n30327 , n17627 , n16095 );
    xnor g30869 ( n24219 , n8924 , n17585 );
    xnor g30870 ( n14582 , n25170 , n19280 );
    not g30871 ( n12215 , n5862 );
    or g30872 ( n18593 , n17619 , n16827 );
    xnor g30873 ( n13982 , n19652 , n23419 );
    xnor g30874 ( n10795 , n22329 , n4982 );
    xnor g30875 ( n16549 , n28059 , n26660 );
    nor g30876 ( n15187 , n13514 , n3870 );
    or g30877 ( n2448 , n6388 , n5120 );
    or g30878 ( n4596 , n15074 , n12778 );
    not g30879 ( n4376 , n17497 );
    or g30880 ( n8226 , n16119 , n5890 );
    not g30881 ( n15762 , n27083 );
    xnor g30882 ( n6259 , n6073 , n25018 );
    xnor g30883 ( n226 , n9043 , n26541 );
    or g30884 ( n7959 , n23342 , n21039 );
    not g30885 ( n15038 , n2444 );
    not g30886 ( n27201 , n15687 );
    xnor g30887 ( n3657 , n7180 , n24578 );
    nor g30888 ( n16723 , n28448 , n14098 );
    and g30889 ( n26995 , n2031 , n30548 );
    xnor g30890 ( n26401 , n31516 , n21229 );
    xnor g30891 ( n20669 , n28828 , n6196 );
    and g30892 ( n2343 , n28373 , n5404 );
    not g30893 ( n17722 , n22664 );
    not g30894 ( n3866 , n3566 );
    not g30895 ( n14030 , n27354 );
    or g30896 ( n23496 , n8019 , n23602 );
    not g30897 ( n4700 , n16119 );
    or g30898 ( n23303 , n26496 , n23802 );
    and g30899 ( n6875 , n29271 , n23763 );
    and g30900 ( n27474 , n2974 , n1259 );
    nor g30901 ( n11934 , n16609 , n21102 );
    or g30902 ( n21477 , n26527 , n11285 );
    or g30903 ( n9249 , n20168 , n1063 );
    nor g30904 ( n17752 , n12037 , n9542 );
    xnor g30905 ( n5102 , n24706 , n21624 );
    not g30906 ( n3762 , n8183 );
    not g30907 ( n30614 , n9455 );
    xor g30908 ( n9929 , n17903 , n16085 );
    xnor g30909 ( n11533 , n24476 , n20116 );
    not g30910 ( n26711 , n24837 );
    and g30911 ( n13077 , n25225 , n21088 );
    xnor g30912 ( n5315 , n20616 , n10269 );
    or g30913 ( n17827 , n14292 , n8894 );
    not g30914 ( n5181 , n17261 );
    or g30915 ( n68 , n20736 , n27037 );
    xnor g30916 ( n30709 , n1742 , n19317 );
    xnor g30917 ( n27639 , n21118 , n15454 );
    or g30918 ( n28677 , n25858 , n8326 );
    xor g30919 ( n11884 , n25824 , n1325 );
    and g30920 ( n7517 , n10402 , n16868 );
    and g30921 ( n5608 , n19556 , n18451 );
    or g30922 ( n9874 , n24942 , n20896 );
    xnor g30923 ( n12797 , n26115 , n11847 );
    xnor g30924 ( n31942 , n593 , n13570 );
    and g30925 ( n20356 , n22954 , n25679 );
    nor g30926 ( n12741 , n6197 , n23857 );
    not g30927 ( n9008 , n3313 );
    xnor g30928 ( n24744 , n24664 , n25134 );
    not g30929 ( n18155 , n15198 );
    or g30930 ( n26156 , n26775 , n1443 );
    and g30931 ( n14399 , n22627 , n22894 );
    not g30932 ( n23202 , n6127 );
    and g30933 ( n16158 , n25209 , n19736 );
    xnor g30934 ( n15509 , n13706 , n871 );
    not g30935 ( n4830 , n8775 );
    not g30936 ( n3967 , n1422 );
    buf g30937 ( n26929 , n9193 );
    and g30938 ( n18315 , n20733 , n11276 );
    xnor g30939 ( n10910 , n17795 , n27493 );
    or g30940 ( n3647 , n4011 , n2619 );
    nor g30941 ( n3028 , n8264 , n15748 );
    or g30942 ( n13007 , n24274 , n7997 );
    xnor g30943 ( n28151 , n25451 , n9966 );
    not g30944 ( n14617 , n24015 );
    or g30945 ( n1589 , n10320 , n16814 );
    xnor g30946 ( n15376 , n16064 , n29014 );
    xnor g30947 ( n9650 , n22378 , n19174 );
    xnor g30948 ( n12895 , n28973 , n7723 );
    and g30949 ( n18218 , n17092 , n17066 );
    nor g30950 ( n6859 , n5995 , n20343 );
    and g30951 ( n28283 , n7039 , n22819 );
    xnor g30952 ( n4324 , n21598 , n1720 );
    not g30953 ( n3244 , n31573 );
    or g30954 ( n15236 , n31913 , n23719 );
    xnor g30955 ( n25657 , n22870 , n891 );
    nor g30956 ( n18407 , n29956 , n9078 );
    xnor g30957 ( n7824 , n28158 , n8014 );
    xnor g30958 ( n31829 , n31759 , n26710 );
    or g30959 ( n25141 , n27782 , n15666 );
    and g30960 ( n25600 , n11555 , n20402 );
    not g30961 ( n8201 , n26684 );
    and g30962 ( n6547 , n9618 , n16341 );
    or g30963 ( n18879 , n21358 , n7338 );
    nor g30964 ( n8882 , n30287 , n19935 );
    or g30965 ( n178 , n18249 , n3344 );
    not g30966 ( n2016 , n16198 );
    and g30967 ( n14845 , n28877 , n12408 );
    or g30968 ( n5171 , n26477 , n8020 );
    nor g30969 ( n2983 , n2615 , n22214 );
    not g30970 ( n3501 , n26191 );
    or g30971 ( n8937 , n1403 , n26979 );
    and g30972 ( n29377 , n6202 , n14232 );
    and g30973 ( n21352 , n28954 , n1596 );
    or g30974 ( n7741 , n7418 , n23580 );
    xor g30975 ( n17052 , n8369 , n28849 );
    xnor g30976 ( n6822 , n30319 , n20391 );
    nor g30977 ( n30093 , n31302 , n31041 );
    not g30978 ( n14661 , n18453 );
    not g30979 ( n20859 , n24669 );
    xnor g30980 ( n7751 , n9210 , n4943 );
    and g30981 ( n29970 , n13142 , n22028 );
    nor g30982 ( n20464 , n20776 , n16889 );
    and g30983 ( n6868 , n18190 , n18950 );
    not g30984 ( n10673 , n23784 );
    and g30985 ( n31316 , n17676 , n113 );
    not g30986 ( n10094 , n24214 );
    not g30987 ( n3569 , n24595 );
    not g30988 ( n30526 , n15759 );
    and g30989 ( n7032 , n1425 , n18199 );
    xnor g30990 ( n31021 , n27889 , n24086 );
    or g30991 ( n20901 , n2087 , n11622 );
    not g30992 ( n11746 , n29499 );
    buf g30993 ( n3787 , n25144 );
    or g30994 ( n7015 , n19999 , n16720 );
    xnor g30995 ( n21968 , n19287 , n22345 );
    xnor g30996 ( n3633 , n30345 , n29089 );
    xnor g30997 ( n7282 , n14048 , n5562 );
    and g30998 ( n19730 , n28760 , n26631 );
    not g30999 ( n30482 , n5610 );
    or g31000 ( n2425 , n26031 , n24480 );
    nor g31001 ( n17871 , n19231 , n27172 );
    and g31002 ( n4868 , n23347 , n30225 );
    nor g31003 ( n24793 , n8724 , n9789 );
    or g31004 ( n4184 , n23053 , n29875 );
    not g31005 ( n7417 , n17165 );
    and g31006 ( n16307 , n31756 , n150 );
    not g31007 ( n29992 , n13923 );
    not g31008 ( n27693 , n16392 );
    not g31009 ( n6482 , n30595 );
    not g31010 ( n20392 , n14610 );
    or g31011 ( n9207 , n13466 , n11235 );
    nor g31012 ( n29880 , n30411 , n15620 );
    and g31013 ( n8664 , n29812 , n15980 );
    not g31014 ( n7596 , n1022 );
    xnor g31015 ( n3331 , n20233 , n7314 );
    nor g31016 ( n25132 , n22858 , n15075 );
    or g31017 ( n999 , n61 , n17919 );
    nor g31018 ( n16374 , n29974 , n14122 );
    nor g31019 ( n18106 , n20236 , n11043 );
    not g31020 ( n26439 , n26966 );
    nor g31021 ( n10283 , n18612 , n21204 );
    or g31022 ( n31071 , n3259 , n13972 );
    xnor g31023 ( n6143 , n14574 , n15914 );
    or g31024 ( n24096 , n19076 , n20817 );
    xnor g31025 ( n3717 , n21933 , n19376 );
    xnor g31026 ( n20251 , n30559 , n16924 );
    nor g31027 ( n23892 , n15948 , n27889 );
    not g31028 ( n14206 , n18413 );
    not g31029 ( n3964 , n7193 );
    not g31030 ( n12613 , n11920 );
    or g31031 ( n7085 , n16411 , n880 );
    or g31032 ( n19136 , n5323 , n30321 );
    not g31033 ( n18356 , n10299 );
    nor g31034 ( n10010 , n11753 , n14606 );
    xnor g31035 ( n948 , n20191 , n20841 );
    not g31036 ( n3696 , n31727 );
    xnor g31037 ( n3185 , n5030 , n9864 );
    or g31038 ( n7063 , n13066 , n9974 );
    xnor g31039 ( n12746 , n27004 , n2067 );
    or g31040 ( n16629 , n11579 , n9760 );
    not g31041 ( n31868 , n12513 );
    not g31042 ( n28629 , n12946 );
    nor g31043 ( n4046 , n16300 , n15401 );
    not g31044 ( n7624 , n10134 );
    xnor g31045 ( n27302 , n20156 , n2898 );
    xor g31046 ( n21383 , n6910 , n9683 );
    nor g31047 ( n26548 , n3416 , n15398 );
    or g31048 ( n18692 , n12501 , n25928 );
    or g31049 ( n24205 , n24958 , n5735 );
    not g31050 ( n13485 , n18984 );
    and g31051 ( n22756 , n30605 , n11103 );
    and g31052 ( n23785 , n14671 , n334 );
    nor g31053 ( n28392 , n16574 , n14619 );
    xnor g31054 ( n6616 , n18279 , n4258 );
    or g31055 ( n27164 , n31290 , n3409 );
    and g31056 ( n1559 , n13922 , n3268 );
    xnor g31057 ( n6784 , n29780 , n18887 );
    not g31058 ( n7858 , n1672 );
    or g31059 ( n19503 , n28445 , n18395 );
    not g31060 ( n28057 , n17221 );
    nor g31061 ( n11119 , n22930 , n23574 );
    not g31062 ( n21815 , n15159 );
    or g31063 ( n985 , n520 , n26270 );
    not g31064 ( n9821 , n26786 );
    not g31065 ( n17364 , n10508 );
    or g31066 ( n18182 , n3810 , n2026 );
    not g31067 ( n16967 , n7687 );
    or g31068 ( n18597 , n6467 , n4717 );
    not g31069 ( n28875 , n18645 );
    not g31070 ( n27927 , n23628 );
    not g31071 ( n22885 , n21735 );
    and g31072 ( n17185 , n29558 , n7700 );
    not g31073 ( n9069 , n4135 );
    and g31074 ( n30234 , n10207 , n14931 );
    xnor g31075 ( n9057 , n7869 , n7808 );
    not g31076 ( n29866 , n17499 );
    not g31077 ( n1796 , n25720 );
    xnor g31078 ( n21793 , n2343 , n14081 );
    and g31079 ( n15225 , n23212 , n3952 );
    xnor g31080 ( n30989 , n31667 , n1587 );
    not g31081 ( n14800 , n5438 );
    or g31082 ( n6116 , n28638 , n6597 );
    not g31083 ( n31514 , n3483 );
    xnor g31084 ( n20424 , n7424 , n10955 );
    xnor g31085 ( n31762 , n3598 , n25150 );
    not g31086 ( n9795 , n9885 );
    xnor g31087 ( n14847 , n14646 , n6717 );
    not g31088 ( n12786 , n14589 );
    and g31089 ( n26503 , n27669 , n25983 );
    nor g31090 ( n1111 , n28610 , n31070 );
    xnor g31091 ( n20775 , n30721 , n771 );
    or g31092 ( n25423 , n20650 , n23371 );
    nor g31093 ( n1014 , n28951 , n2629 );
    or g31094 ( n23837 , n22571 , n15852 );
    xnor g31095 ( n31182 , n4699 , n17367 );
    xnor g31096 ( n21262 , n15178 , n7701 );
    xnor g31097 ( n22874 , n10622 , n21973 );
    not g31098 ( n5249 , n27907 );
    and g31099 ( n5413 , n23654 , n7370 );
    xnor g31100 ( n31170 , n14524 , n9414 );
    or g31101 ( n8438 , n823 , n7998 );
    xnor g31102 ( n2408 , n26230 , n30359 );
    xor g31103 ( n6510 , n13703 , n20 );
    or g31104 ( n21423 , n27153 , n3338 );
    xnor g31105 ( n27033 , n28489 , n2386 );
    not g31106 ( n4854 , n15435 );
    or g31107 ( n17449 , n26261 , n16540 );
    or g31108 ( n14863 , n19930 , n19553 );
    not g31109 ( n21279 , n6358 );
    xnor g31110 ( n30423 , n26583 , n7304 );
    not g31111 ( n22553 , n9826 );
    and g31112 ( n23339 , n15034 , n16399 );
    not g31113 ( n17469 , n6128 );
    not g31114 ( n4970 , n19558 );
    xnor g31115 ( n19981 , n6428 , n11028 );
    or g31116 ( n6073 , n21692 , n24555 );
    xnor g31117 ( n19361 , n23419 , n8867 );
    or g31118 ( n12046 , n8547 , n829 );
    or g31119 ( n8389 , n6142 , n20802 );
    or g31120 ( n9560 , n2636 , n19209 );
    xnor g31121 ( n28948 , n2541 , n9371 );
    or g31122 ( n15913 , n812 , n11028 );
    xnor g31123 ( n17251 , n7434 , n3106 );
    not g31124 ( n9956 , n8479 );
    not g31125 ( n26489 , n6972 );
    xnor g31126 ( n6826 , n24469 , n15449 );
    or g31127 ( n781 , n21930 , n28221 );
    not g31128 ( n27460 , n5638 );
    or g31129 ( n1884 , n2510 , n16299 );
    and g31130 ( n28639 , n361 , n22852 );
    and g31131 ( n6269 , n4436 , n15709 );
    not g31132 ( n22816 , n29183 );
    xnor g31133 ( n8826 , n17931 , n28898 );
    xnor g31134 ( n20089 , n31781 , n16790 );
    and g31135 ( n17567 , n3898 , n11708 );
    not g31136 ( n21232 , n24873 );
    nor g31137 ( n7727 , n20388 , n29131 );
    not g31138 ( n19010 , n9710 );
    nor g31139 ( n12928 , n20427 , n6078 );
    not g31140 ( n2853 , n25164 );
    not g31141 ( n26300 , n22227 );
    not g31142 ( n11438 , n12777 );
    buf g31143 ( n2515 , n3261 );
    nor g31144 ( n15377 , n22875 , n25688 );
    or g31145 ( n29232 , n19003 , n23398 );
    nor g31146 ( n26412 , n21216 , n18924 );
    xnor g31147 ( n11333 , n20262 , n26961 );
    and g31148 ( n11766 , n27060 , n30734 );
    not g31149 ( n9639 , n22968 );
    or g31150 ( n12008 , n16113 , n2842 );
    or g31151 ( n22476 , n31725 , n21941 );
    and g31152 ( n21318 , n18220 , n14818 );
    and g31153 ( n4456 , n6287 , n4065 );
    xnor g31154 ( n9217 , n10843 , n3622 );
    not g31155 ( n287 , n1166 );
    or g31156 ( n15532 , n20062 , n19192 );
    not g31157 ( n31856 , n20442 );
    or g31158 ( n15938 , n28856 , n3268 );
    or g31159 ( n1572 , n10664 , n29285 );
    xnor g31160 ( n12751 , n24246 , n11574 );
    or g31161 ( n7041 , n14976 , n19778 );
    or g31162 ( n17404 , n20367 , n8855 );
    or g31163 ( n18183 , n16084 , n29201 );
    xnor g31164 ( n14658 , n12558 , n27453 );
    or g31165 ( n3876 , n17843 , n9179 );
    xnor g31166 ( n14398 , n24354 , n30010 );
    xnor g31167 ( n11852 , n23973 , n27433 );
    and g31168 ( n14088 , n16959 , n7316 );
    xnor g31169 ( n4196 , n6455 , n20210 );
    nor g31170 ( n16489 , n2934 , n16342 );
    and g31171 ( n21637 , n5520 , n4800 );
    xor g31172 ( n3079 , n2870 , n2934 );
    or g31173 ( n21792 , n28565 , n3796 );
    xnor g31174 ( n10226 , n27445 , n2424 );
    not g31175 ( n407 , n14705 );
    not g31176 ( n4567 , n8908 );
    and g31177 ( n17245 , n23033 , n26649 );
    not g31178 ( n7353 , n21760 );
    not g31179 ( n19545 , n14901 );
    xnor g31180 ( n20444 , n31257 , n11016 );
    not g31181 ( n24111 , n11837 );
    not g31182 ( n16525 , n20736 );
    and g31183 ( n17283 , n7304 , n12048 );
    and g31184 ( n23875 , n19722 , n23619 );
    not g31185 ( n15414 , n4570 );
    and g31186 ( n27599 , n31838 , n28692 );
    xnor g31187 ( n16269 , n19714 , n14129 );
    xnor g31188 ( n28178 , n19734 , n9358 );
    or g31189 ( n30054 , n25123 , n24075 );
    not g31190 ( n3963 , n6320 );
    not g31191 ( n8701 , n24442 );
    and g31192 ( n15246 , n22068 , n26693 );
    not g31193 ( n28008 , n24524 );
    and g31194 ( n18526 , n13341 , n12103 );
endmodule
